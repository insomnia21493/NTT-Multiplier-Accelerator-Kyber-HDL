library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ROM is
port (
    clk   : in std_logic;
    addr  : in std_logic_vector(7 downto 0);
    dout  : out std_logic_vector(11 downto 0)
);
end ROM;



architecture RTL of ROM is
    type MEMORY is array (0 to 255) of std_logic_vector(11 downto 0);
    constant ROM_mem : MEMORY := (
		x"674",
		x"6c1",
		x"a14",
		x"cd9",
		x"a52",
		x"276",
		x"769",
		x"350",
		x"426",
		x"77f",
		x"0c1",
		x"31d",
		x"ae2",
		x"cbc",
		x"239",
		x"6d2",
		x"128",
		x"98f",
		x"53b",
		x"5c4",
		x"be6",
		x"038",
		x"8c0",
		x"535",
		x"592",
		x"82e",
		x"217",
		x"b42",
		x"959",
		x"b3f",
		x"7b6",
		x"335",
		x"121",
		x"14b",
		x"cb5",
		x"6dc",
		x"4ad",
		x"900",
		x"8e5",
		x"807",
		x"28a",
		x"7b9",
		x"9d1",
		x"278",
		x"b31",
		x"021",
		x"528",
		x"77b",
		x"90f",
		x"59b",
		x"327",
		x"1c4",
		x"59e",
		x"b34",
		x"5fe",
		x"962",
		x"a57",
		x"a39",
		x"5c9",
		x"288",
		x"9aa",
		x"c26",
		x"4cb",
		x"38e",
		x"011",
		x"ac9",
		x"247",
		x"a59",
		x"665",
		x"2d3",
		x"8f0",
		x"44c",
		x"581",
		x"a66",
		x"cd1",
		x"0e9",
		x"2f4",
		x"86c",
		x"bc7",
		x"bea",
		x"6a7",
		x"673",
		x"ae5",
		x"6fd",
		x"737",
		x"3b8",
		x"5b5",
		x"a7f",
		x"3ab",
		x"904",
		x"985",
		x"954",
		x"2dd",
		x"921",
		x"10c",
		x"281",
		x"630",
		x"8fa",
		x"7f5",
		x"c94",
		x"177",
		x"9f5",
		x"82a",
		x"66d",
		x"427",
		x"13f",
		x"ad5",
		x"2f5",
		x"833",
		x"231",
		x"9a2",
		x"a22",
		x"af4",
		x"444",
		x"193",
		x"402",
		x"477",
		x"866",
		x"ad7",
		x"376",
		x"6ba",
		x"4bc",
		x"752",
		x"405",
		x"83e",
		x"b77",
		x"375",
		x"86a",
-- rest is negative zetas		
		x"ce7",
		x"640",
		x"2ed",
		x"028",
		x"2af",
		x"a8b",
		x"598",
		x"9b1",
		x"8db",
		x"582",
		x"c40",
		x"9e4",
		x"21f",
		x"045",
		x"ac8",
		x"62f",
		x"bd9",
		x"372",
		x"7c6",
		x"73d",
		x"11b",
		x"cc9",
		x"441",
		x"7cc",
		x"76f",
		x"4d3",
		x"aea",
		x"1bf",
		x"3a8",
		x"1c2",
		x"54b",
		x"9cc",
		x"be0",
		x"bb6",
		x"04c",
		x"625",
		x"854",
		x"401",
		x"41c",
		x"4fa",
		x"a77",
		x"548",
		x"330",
		x"a89",
		x"1d0",
		x"ce0",
		x"7d9",
		x"586",
		x"3f2",
		x"766",
		x"9da",
		x"b3d",
		x"763",
		x"1cd",
		x"703",
		x"39f",
		x"2aa",
		x"2c8",
		x"738",
		x"a79",
		x"357",
		x"0db",
		x"836",
		x"973",
		x"cf0",
		x"238",
		x"aba",
		x"2a8",
		x"69c",
		x"a2e",
		x"411",
		x"8b5",
		x"780",
		x"29b",
		x"030",
		x"c18",
		x"a0d",
		x"495",
		x"13a",
		x"117",
		x"65a",
		x"68e",
		x"21c",
		x"604",
		x"5ca",
		x"949",
		x"74c",
		x"282",
		x"956",
		x"3fd",
		x"37c",
		x"3ad",
		x"a24",
		x"3e0",
		x"bf5",
		x"a80",
		x"6d1",
		x"407",
		x"50c",
		x"06d",
		x"b8a",
		x"30c",
		x"4d7",
		x"694",
		x"8da",
		x"bc2",
		x"22c",
		x"a0c",
		x"4ce",
		x"ad0",
		x"35f",
		x"2df",
		x"20d",
		x"8bd",
		x"b6e",
		x"8ff",
		x"88a",
		x"49b",
		x"22a",
		x"98b",
		x"647",
		x"845",
		x"5af",
		x"8fc",
		x"4c3",
		x"18a",
		x"98c",
		x"497"	

    );
begin
    process(clk)
		begin
			if(clk'event and clk='1') then
				dout <= ROM_mem(conv_integer(addr));
			end if;
		end process;

end architecture RTL;