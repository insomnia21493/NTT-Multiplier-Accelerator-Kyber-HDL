LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL; 
LIBRARY work;
USE work.ALL;


ENTITY ntttb IS END ntttb;



ARCHITECTURE test OF ntttb IS

    COMPONENT ntt IS
			PORT(
				clk         	:   IN  	std_logic;
				nrst        	:   IN  	std_logic;
				en	        	:   IN  	std_logic;
				mode	        :	IN		std_logic_vector(1 downto 0);
				WE				:	IN		std_logic;
				Address			:	IN		std_logic_vector(8 downto 0);
				Data_In			:	IN		std_logic_vector(11 downto 0);  
				Data_Out		:	OUT		std_logic_vector(11 downto 0);				
				busy        	:   OUT 	std_logic;
				done        	:   OUT 	std_logic
				
				
				);

		END COMPONENT;
	
	

	
	SIGNAL	tbclk       	:   std_logic:='1';
	SIGNAL	tbnrst      	:   std_logic;
	SIGNAL	tben	        	:  	std_logic;
	SIGNAL	tbmode	        :	std_logic_vector(1 downto 0);
	SIGNAL	tbWE			:	std_logic;
	SIGNAL	tbAddress		:	std_logic_vector(8 downto 0);
	SIGNAL	tbData_In		:	std_logic_vector(11 downto 0);  
	SIGNAL	tbData_Out		:	std_logic_vector(11 downto 0);		
	SIGNAL  tbbusy        	:  	std_logic;
	SIGNAL  tbdone        	:  	std_logic;
	
	
	
BEGIN  
  
  	ntt_for_test: ntt PORT MAP (
							
							clk      => tbclk	  ,     
							nrst     => tbnrst    ,
							en	     => tben	  ,
							mode	 => tbmode	  ,
							WE		 => tbWE	  ,
							Address	 => tbAddress ,
							Data_In	 => tbData_In ,
							Data_Out => tbData_Out,
							busy     => tbbusy    ,
							done     => tbdone    
														
							);
	


  tbclk <= NOT tbclk AFTER 5 ns;

PROCESS
	BEGIN
	
		
		tbnrst <= '0';

	wait for 10 ns;
		
		tbnrst <= '1';
		
		tbmode	<="00";
	
	wait for 10 ns;
	
		

		tbData_In  <="110000111101";
		tbAddress  <="000000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000101001";
		tbAddress  <="000000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000010101";
		tbAddress  <="000000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110111101";
		tbAddress  <="000000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010011111";
		tbAddress  <="000000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001001111";
		tbAddress  <="000000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010001101";
		tbAddress  <="000000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000010110";
		tbAddress  <="000000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010101100";
		tbAddress  <="000001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110100101";
		tbAddress  <="000001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011100100";
		tbAddress  <="000001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101101101";
		tbAddress  <="000001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111000110";
		tbAddress  <="000001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111110100";
		tbAddress  <="000001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001111001";
		tbAddress  <="000001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000100111";
		tbAddress  <="000001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100000";
		tbAddress  <="000010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011010101";
		tbAddress  <="000010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100100101";
		tbAddress  <="000010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011001001";
		tbAddress  <="000010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000000010";
		tbAddress  <="000010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100111100";
		tbAddress  <="000010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011011101";
		tbAddress  <="000010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110011101";
		tbAddress  <="000010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010101000";
		tbAddress  <="000011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001000100";
		tbAddress  <="000011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110001011";
		tbAddress  <="000011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100111";
		tbAddress  <="000011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100111001";
		tbAddress  <="000011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011100011";
		tbAddress  <="000011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011001001";
		tbAddress  <="000011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001001110";
		tbAddress  <="000011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100001100";
		tbAddress  <="000100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011100110";
		tbAddress  <="000100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010001010";
		tbAddress  <="000100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001000001";
		tbAddress  <="000100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001100001";
		tbAddress  <="000100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100010010";
		tbAddress  <="000100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000010111";
		tbAddress  <="000100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000101010";
		tbAddress  <="000100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100110010";
		tbAddress  <="000101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101011001";
		tbAddress  <="000101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011000011";
		tbAddress  <="000101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010101100";
		tbAddress  <="000101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001000000";
		tbAddress  <="000101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000011011";
		tbAddress  <="000101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111011011";
		tbAddress  <="000101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100101101";
		tbAddress  <="000101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010010110";
		tbAddress  <="000110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010110001";
		tbAddress  <="000110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010100";
		tbAddress  <="000110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101111101";
		tbAddress  <="000110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110111000";
		tbAddress  <="000110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110110110";
		tbAddress  <="000110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110001011";
		tbAddress  <="000110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101101011";
		tbAddress  <="000110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000110011";
		tbAddress  <="000111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110011000";
		tbAddress  <="000111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010011";
		tbAddress  <="000111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010101001";
		tbAddress  <="000111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111101111";
		tbAddress  <="000111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011010001";
		tbAddress  <="000111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110001111";
		tbAddress  <="000111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011110100";
		tbAddress  <="000111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010010";
		tbAddress  <="001000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100001100";
		tbAddress  <="001000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010011000";
		tbAddress  <="001000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011010011";
		tbAddress  <="001000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010100000";
		tbAddress  <="001000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100001";
		tbAddress  <="001000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000101110";
		tbAddress  <="001000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011011011";
		tbAddress  <="001000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101101000";
		tbAddress  <="001001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111000111";
		tbAddress  <="001001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100000001";
		tbAddress  <="001001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101001110";
		tbAddress  <="001001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101110110";
		tbAddress  <="001001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111010101";
		tbAddress  <="001001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110000";
		tbAddress  <="001001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010111110";
		tbAddress  <="001001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001010001";
		tbAddress  <="001010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001010110";
		tbAddress  <="001010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001101000";
		tbAddress  <="001010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101110001";
		tbAddress  <="001010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111010100";
		tbAddress  <="001010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101000100";
		tbAddress  <="001010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110100110";
		tbAddress  <="001010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001001110";
		tbAddress  <="001010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010011111";
		tbAddress  <="001011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100110100";
		tbAddress  <="001011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011000011";
		tbAddress  <="001011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011111010";
		tbAddress  <="001011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010000110";
		tbAddress  <="001011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010010101";
		tbAddress  <="001011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110010111";
		tbAddress  <="001011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010100111";
		tbAddress  <="001011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010110010";
		tbAddress  <="001100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001111001";
		tbAddress  <="001100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101110111";
		tbAddress  <="001100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010110101";
		tbAddress  <="001100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000111111";
		tbAddress  <="001100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100101001";
		tbAddress  <="001100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110110110";
		tbAddress  <="001100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100100101";
		tbAddress  <="001100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000011101";
		tbAddress  <="001101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110101010";
		tbAddress  <="001101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000001100";
		tbAddress  <="001101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110011110";
		tbAddress  <="001101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010000111";
		tbAddress  <="001101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001010001";
		tbAddress  <="001101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011000110";
		tbAddress  <="001101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000011001";
		tbAddress  <="001101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110011111";
		tbAddress  <="001110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111000000";
		tbAddress  <="001110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110110";
		tbAddress  <="001110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011011011";
		tbAddress  <="001110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010000101";
		tbAddress  <="001110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001001010";
		tbAddress  <="001110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100001011";
		tbAddress  <="001110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001110001";
		tbAddress  <="001110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110111001";
		tbAddress  <="001111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110111001";
		tbAddress  <="001111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101001011";
		tbAddress  <="001111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000111101";
		tbAddress  <="001111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000000100";
		tbAddress  <="001111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111101100";
		tbAddress  <="001111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110101100";
		tbAddress  <="001111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111110110";
		tbAddress  <="001111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010110011";
		tbAddress  <="010000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110010110";
		tbAddress  <="010000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001101100";
		tbAddress  <="010000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111111010";
		tbAddress  <="010000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111111100";
		tbAddress  <="010000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100100110";
		tbAddress  <="010000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011011010";
		tbAddress  <="010000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010000110";
		tbAddress  <="010000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001111111";
		tbAddress  <="010001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001011111";
		tbAddress  <="010001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001000011";
		tbAddress  <="010001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100111011";
		tbAddress  <="010001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001100110";
		tbAddress  <="010001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010100110";
		tbAddress  <="010001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111001001";
		tbAddress  <="010001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111001110";
		tbAddress  <="010001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111000101";
		tbAddress  <="010010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110001101";
		tbAddress  <="010010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010010111";
		tbAddress  <="010010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001010100";
		tbAddress  <="010010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010101100";
		tbAddress  <="010010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000000001";
		tbAddress  <="010010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011011111";
		tbAddress  <="010010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001010100";
		tbAddress  <="010010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000001110";
		tbAddress  <="010011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010010000";
		tbAddress  <="010011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000110011";
		tbAddress  <="010011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000011101";
		tbAddress  <="010011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000111010";
		tbAddress  <="010011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010001000";
		tbAddress  <="010011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101100011";
		tbAddress  <="010011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000110011";
		tbAddress  <="010011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010110110";
		tbAddress  <="010100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111100100";
		tbAddress  <="010100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010001011";
		tbAddress  <="010100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011101010";
		tbAddress  <="010100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100001";
		tbAddress  <="010100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100001";
		tbAddress  <="010100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010110110";
		tbAddress  <="010100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000111001";
		tbAddress  <="010100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101010101";
		tbAddress  <="010101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110000101";
		tbAddress  <="010101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000001101";
		tbAddress  <="010101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001000111";
		tbAddress  <="010101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001010011";
		tbAddress  <="010101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010110";
		tbAddress  <="010101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100001011";
		tbAddress  <="010101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011001000";
		tbAddress  <="010101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001000110";
		tbAddress  <="010110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000000110";
		tbAddress  <="010110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110111111";
		tbAddress  <="010110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011000110";
		tbAddress  <="010110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011000101";
		tbAddress  <="010110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010010";
		tbAddress  <="010110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111111001";
		tbAddress  <="010110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110101010";
		tbAddress  <="010110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010100110";
		tbAddress  <="010111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111110011";
		tbAddress  <="010111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011101110";
		tbAddress  <="010111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111011100";
		tbAddress  <="010111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000010010";
		tbAddress  <="010111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000100001";
		tbAddress  <="010111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100010000";
		tbAddress  <="010111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111111010";
		tbAddress  <="010111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011100110";
		tbAddress  <="011000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100001000";
		tbAddress  <="011000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101011000";
		tbAddress  <="011000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101110101";
		tbAddress  <="011000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101000110";
		tbAddress  <="011000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000101100";
		tbAddress  <="011000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101011001";
		tbAddress  <="011000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100010000";
		tbAddress  <="011000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001110011";
		tbAddress  <="011001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000000101";
		tbAddress  <="011001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000001011";
		tbAddress  <="011001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001100110";
		tbAddress  <="011001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101001110";
		tbAddress  <="011001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111011001";
		tbAddress  <="011001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000001110";
		tbAddress  <="011001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100000001";
		tbAddress  <="011001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100100000";
		tbAddress  <="011010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111010011";
		tbAddress  <="011010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100001001";
		tbAddress  <="011010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010110000";
		tbAddress  <="011010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000011111";
		tbAddress  <="011010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010011011";
		tbAddress  <="011010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001001100";
		tbAddress  <="011010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011011010";
		tbAddress  <="011010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010110110";
		tbAddress  <="011011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011100001";
		tbAddress  <="011011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010011110";
		tbAddress  <="011011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001001111";
		tbAddress  <="011011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011001011";
		tbAddress  <="011011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111001010";
		tbAddress  <="011011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011001010";
		tbAddress  <="011011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001110010";
		tbAddress  <="011011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001001110";
		tbAddress  <="011100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010110010";
		tbAddress  <="011100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101100101";
		tbAddress  <="011100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001010010";
		tbAddress  <="011100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100111010";
		tbAddress  <="011100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001000111";
		tbAddress  <="011100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101100000";
		tbAddress  <="011100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101011101";
		tbAddress  <="011100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100010110";
		tbAddress  <="011101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000111111";
		tbAddress  <="011101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100100001";
		tbAddress  <="011101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000001001";
		tbAddress  <="011101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100111011";
		tbAddress  <="011101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111110";
		tbAddress  <="011101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010111111";
		tbAddress  <="011101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011001010";
		tbAddress  <="011101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001011001";
		tbAddress  <="011110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101001111";
		tbAddress  <="011110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011010110";
		tbAddress  <="011110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011111011";
		tbAddress  <="011110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100101010";
		tbAddress  <="011110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100011110";
		tbAddress  <="011110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100001001";
		tbAddress  <="011110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111110000";
		tbAddress  <="011110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001000001";
		tbAddress  <="011111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100100101";
		tbAddress  <="011111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100110001";
		tbAddress  <="011111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111000";
		tbAddress  <="011111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100011110";
		tbAddress  <="011111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000100101";
		tbAddress  <="011111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010010111";
		tbAddress  <="011111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001011001";
		tbAddress  <="011111111";
		tbWE  <='1';
		wait for 10 ns;	
		tbWE  <='0';
		tbmode <= "00";
		tben<='1';
		
		wait for 10 ns;	
		
		tben<='0';
		
		wait for 20000 ns;	
		
		tbmode <= "10";
		tben<='1';
		
		wait for 10 ns;	
		
		tben<='1';
		
		
		wait for 10 ns;	
		
		tben<='0';
		
		wait for 20000 ns;	
		
		
		
		tbData_In  <="101011110000";
		tbAddress  <="000000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001010010";
		tbAddress  <="000000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101001110";
		tbAddress  <="000000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000010001";
		tbAddress  <="000000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110110";
		tbAddress  <="000000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011110000";
		tbAddress  <="000000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101110101";
		tbAddress  <="000000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011111010";
		tbAddress  <="000000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001111010";
		tbAddress  <="000001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011110111";
		tbAddress  <="000001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110000100";
		tbAddress  <="000001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110101100";
		tbAddress  <="000001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111110010";
		tbAddress  <="000001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100101101";
		tbAddress  <="000001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011010111";
		tbAddress  <="000001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101110110";
		tbAddress  <="000001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010101010";
		tbAddress  <="000010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001001010";
		tbAddress  <="000010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000110000";
		tbAddress  <="000010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111001110";
		tbAddress  <="000010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101000110";
		tbAddress  <="000010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011000110";
		tbAddress  <="000010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010000001";
		tbAddress  <="000010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000011111";
		tbAddress  <="000010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111111010";
		tbAddress  <="000011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111011011";
		tbAddress  <="000011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101111011";
		tbAddress  <="000011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101100101";
		tbAddress  <="000011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100001001";
		tbAddress  <="000011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100111000";
		tbAddress  <="000011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011100001";
		tbAddress  <="000011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111001000";
		tbAddress  <="000011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101111101";
		tbAddress  <="000100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111001000";
		tbAddress  <="000100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011011001";
		tbAddress  <="000100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111010111";
		tbAddress  <="000100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111000101";
		tbAddress  <="000100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011110111";
		tbAddress  <="000100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111001101";
		tbAddress  <="000100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010000000";
		tbAddress  <="000100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001000101";
		tbAddress  <="000101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001011010";
		tbAddress  <="000101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111101000";
		tbAddress  <="000101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010100000";
		tbAddress  <="000101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000010000";
		tbAddress  <="000101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101011010";
		tbAddress  <="000101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000001100";
		tbAddress  <="000101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001001000";
		tbAddress  <="000101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011000100";
		tbAddress  <="000110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111101000";
		tbAddress  <="000110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110001001";
		tbAddress  <="000110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010010001";
		tbAddress  <="000110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100110111";
		tbAddress  <="000110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011010001";
		tbAddress  <="000110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010110";
		tbAddress  <="000110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001100100";
		tbAddress  <="000110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110110011";
		tbAddress  <="000111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001010000";
		tbAddress  <="000111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001000101";
		tbAddress  <="000111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111100001";
		tbAddress  <="000111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001011010";
		tbAddress  <="000111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100110001";
		tbAddress  <="000111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101001100";
		tbAddress  <="000111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100110100";
		tbAddress  <="000111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110100101";
		tbAddress  <="001000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110111110";
		tbAddress  <="001000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011111010";
		tbAddress  <="001000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001100100";
		tbAddress  <="001000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001011110";
		tbAddress  <="001000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110010010";
		tbAddress  <="001000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000110001";
		tbAddress  <="001000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010011110";
		tbAddress  <="001000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011011001";
		tbAddress  <="001001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011010011";
		tbAddress  <="001001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100001111";
		tbAddress  <="001001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111001010";
		tbAddress  <="001001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001100000";
		tbAddress  <="001001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010010001";
		tbAddress  <="001001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000000101";
		tbAddress  <="001001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001110111";
		tbAddress  <="001001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100000";
		tbAddress  <="001010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011000000";
		tbAddress  <="001010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000011000";
		tbAddress  <="001010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101110110";
		tbAddress  <="001010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111000111";
		tbAddress  <="001010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100111000";
		tbAddress  <="001010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111111100";
		tbAddress  <="001010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100000001";
		tbAddress  <="001010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100110001";
		tbAddress  <="001011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111100110";
		tbAddress  <="001011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110011011";
		tbAddress  <="001011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101111000";
		tbAddress  <="001011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010101011";
		tbAddress  <="001011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100001100";
		tbAddress  <="001011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111101101";
		tbAddress  <="001011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001000110";
		tbAddress  <="001011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001100011";
		tbAddress  <="001100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000001010";
		tbAddress  <="001100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010000010";
		tbAddress  <="001100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110000001";
		tbAddress  <="001100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001101101";
		tbAddress  <="001100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010000010";
		tbAddress  <="001100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101000010";
		tbAddress  <="001100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000111110";
		tbAddress  <="001100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011110111";
		tbAddress  <="001101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001000100";
		tbAddress  <="001101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111101000";
		tbAddress  <="001101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100011011";
		tbAddress  <="001101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001110001";
		tbAddress  <="001101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011010101";
		tbAddress  <="001101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000011010";
		tbAddress  <="001101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010111010";
		tbAddress  <="001101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000101011";
		tbAddress  <="001110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110101000";
		tbAddress  <="001110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000110111";
		tbAddress  <="001110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111010101";
		tbAddress  <="001110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111100011";
		tbAddress  <="001110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001101111";
		tbAddress  <="001110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101100001";
		tbAddress  <="001110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000110110";
		tbAddress  <="001110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100010";
		tbAddress  <="001111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100101";
		tbAddress  <="001111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000011011";
		tbAddress  <="001111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101110011";
		tbAddress  <="001111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011001110";
		tbAddress  <="001111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000100010";
		tbAddress  <="001111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010011011";
		tbAddress  <="001111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000100001";
		tbAddress  <="001111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010101111";
		tbAddress  <="010000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001010011";
		tbAddress  <="010000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111111001";
		tbAddress  <="010000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001100000";
		tbAddress  <="010000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001111011";
		tbAddress  <="010000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101001011";
		tbAddress  <="010000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011111011";
		tbAddress  <="010000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000100000";
		tbAddress  <="010000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111101000";
		tbAddress  <="010001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010101010";
		tbAddress  <="010001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101111110";
		tbAddress  <="010001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000010010";
		tbAddress  <="010001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001010101";
		tbAddress  <="010001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010110101";
		tbAddress  <="010001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100111011";
		tbAddress  <="010001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000000110";
		tbAddress  <="010001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100001111";
		tbAddress  <="010010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100110011";
		tbAddress  <="010010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010110011";
		tbAddress  <="010010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010111111";
		tbAddress  <="010010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111000001";
		tbAddress  <="010010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011110101";
		tbAddress  <="010010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110000100";
		tbAddress  <="010010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100110011";
		tbAddress  <="010010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001001001";
		tbAddress  <="010011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001110001";
		tbAddress  <="010011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010111111";
		tbAddress  <="010011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101101110";
		tbAddress  <="010011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110001110";
		tbAddress  <="010011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001111100";
		tbAddress  <="010011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101110000";
		tbAddress  <="010011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000011101";
		tbAddress  <="010011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000101000";
		tbAddress  <="010100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101001101";
		tbAddress  <="010100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101011100";
		tbAddress  <="010100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110010100";
		tbAddress  <="010100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001010011";
		tbAddress  <="010100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111100011";
		tbAddress  <="010100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101001111";
		tbAddress  <="010100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100100110";
		tbAddress  <="010100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011101111";
		tbAddress  <="010101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010000100";
		tbAddress  <="010101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100101100";
		tbAddress  <="010101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000110011";
		tbAddress  <="010101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000101001";
		tbAddress  <="010101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101001000";
		tbAddress  <="010101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111110010";
		tbAddress  <="010101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010110101";
		tbAddress  <="010101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111001010";
		tbAddress  <="010110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001101000";
		tbAddress  <="010110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100100001";
		tbAddress  <="010110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110111110";
		tbAddress  <="010110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010110100";
		tbAddress  <="010110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100000010";
		tbAddress  <="010110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111011010";
		tbAddress  <="010110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100110100";
		tbAddress  <="010110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001111001";
		tbAddress  <="010111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100000100";
		tbAddress  <="010111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110110111";
		tbAddress  <="010111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111000010";
		tbAddress  <="010111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110001011";
		tbAddress  <="010111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110110010";
		tbAddress  <="010111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110110000";
		tbAddress  <="010111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010000100";
		tbAddress  <="010111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011100110";
		tbAddress  <="011000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101000000";
		tbAddress  <="011000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111000";
		tbAddress  <="011000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011111011";
		tbAddress  <="011000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001001110";
		tbAddress  <="011000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011010110";
		tbAddress  <="011000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010000011";
		tbAddress  <="011000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011101100";
		tbAddress  <="011000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001111001";
		tbAddress  <="011001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110101000";
		tbAddress  <="011001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001001001";
		tbAddress  <="011001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110011000";
		tbAddress  <="011001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101011001";
		tbAddress  <="011001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111111010";
		tbAddress  <="011001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111010100";
		tbAddress  <="011001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011011110";
		tbAddress  <="011001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000011000";
		tbAddress  <="011010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011110011";
		tbAddress  <="011010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100101010";
		tbAddress  <="011010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111111110";
		tbAddress  <="011010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111000001";
		tbAddress  <="011010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011000110";
		tbAddress  <="011010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110110100";
		tbAddress  <="011010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011110000";
		tbAddress  <="011010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000010101";
		tbAddress  <="011011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001011001";
		tbAddress  <="011011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011011110";
		tbAddress  <="011011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011110000";
		tbAddress  <="011011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101100110";
		tbAddress  <="011011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111110101";
		tbAddress  <="011011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101011000";
		tbAddress  <="011011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001010011";
		tbAddress  <="011011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011011000";
		tbAddress  <="011100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011101001";
		tbAddress  <="011100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011100001";
		tbAddress  <="011100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011110000";
		tbAddress  <="011100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111110000";
		tbAddress  <="011100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010101100";
		tbAddress  <="011100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000011100";
		tbAddress  <="011100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011001101";
		tbAddress  <="011100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010111010";
		tbAddress  <="011101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010001000";
		tbAddress  <="011101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110001100";
		tbAddress  <="011101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000101000";
		tbAddress  <="011101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010111000";
		tbAddress  <="011101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100000000";
		tbAddress  <="011101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010101100";
		tbAddress  <="011101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000100100";
		tbAddress  <="011101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001010011";
		tbAddress  <="011110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001001000";
		tbAddress  <="011110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101110000";
		tbAddress  <="011110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101000010";
		tbAddress  <="011110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100111101";
		tbAddress  <="011110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101101101";
		tbAddress  <="011110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110111";
		tbAddress  <="011110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111011010";
		tbAddress  <="011110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100001010111";
		tbAddress  <="011111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010000010";
		tbAddress  <="011111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110000100";
		tbAddress  <="011111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100000000";
		tbAddress  <="011111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101001010";
		tbAddress  <="011111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010110000";
		tbAddress  <="011111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110010110";
		tbAddress  <="011111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111101110";
		tbAddress  <="011111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101100110";
		tbAddress  <="100000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010011001";
		tbAddress  <="100000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111101000";
		tbAddress  <="100000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111010001";
		tbAddress  <="100000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100011000";
		tbAddress  <="100000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011100110";
		tbAddress  <="100000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011111000";
		tbAddress  <="100000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110100111";
		tbAddress  <="100000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011100001";
		tbAddress  <="100001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010101010";
		tbAddress  <="100001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010001101";
		tbAddress  <="100001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110010110";
		tbAddress  <="100001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101100111";
		tbAddress  <="100001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110110100";
		tbAddress  <="100001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111100001";
		tbAddress  <="100001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011111110";
		tbAddress  <="100001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001010011";
		tbAddress  <="100010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001111111";
		tbAddress  <="100010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010101110";
		tbAddress  <="100010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100110";
		tbAddress  <="100010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101011111";
		tbAddress  <="100010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111111101";
		tbAddress  <="100010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110000110";
		tbAddress  <="100010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111011001";
		tbAddress  <="100010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110011100";
		tbAddress  <="100011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110000110";
		tbAddress  <="100011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011001100";
		tbAddress  <="100011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011001001";
		tbAddress  <="100011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111001000";
		tbAddress  <="100011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010000011";
		tbAddress  <="100011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010011000";
		tbAddress  <="100011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000001110";
		tbAddress  <="100011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011011101";
		tbAddress  <="100100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101000011";
		tbAddress  <="100100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000000000";
		tbAddress  <="100100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011101100";
		tbAddress  <="100100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010111100";
		tbAddress  <="100100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010010111";
		tbAddress  <="100100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001011010";
		tbAddress  <="100100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001011110";
		tbAddress  <="100100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100100110";
		tbAddress  <="100101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111101110";
		tbAddress  <="100101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001110000";
		tbAddress  <="100101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010110000";
		tbAddress  <="100101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000010010";
		tbAddress  <="100101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011000110";
		tbAddress  <="100101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111011011";
		tbAddress  <="100101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010110010";
		tbAddress  <="100101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111010001";
		tbAddress  <="100110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011010111";
		tbAddress  <="100110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001000100";
		tbAddress  <="100110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011000000";
		tbAddress  <="100110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111000010";
		tbAddress  <="100110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001000100100";
		tbAddress  <="100110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110000011";
		tbAddress  <="100110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111011011";
		tbAddress  <="100110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110101001";
		tbAddress  <="100111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001100010";
		tbAddress  <="100111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110100100";
		tbAddress  <="100111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001111010011";
		tbAddress  <="100111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000101001";
		tbAddress  <="100111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011111001";
		tbAddress  <="100111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011100111";
		tbAddress  <="100111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011101101101";
		tbAddress  <="100111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011001110";
		tbAddress  <="101000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110011111";
		tbAddress  <="101000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000011011";
		tbAddress  <="101000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011101001";
		tbAddress  <="101000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001011000";
		tbAddress  <="101000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010100001";
		tbAddress  <="101000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101100011";
		tbAddress  <="101000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000010101";
		tbAddress  <="101000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001110011";
		tbAddress  <="101001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010010011";
		tbAddress  <="101001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000101000";
		tbAddress  <="101001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111110100";
		tbAddress  <="101001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101111111";
		tbAddress  <="101001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011000111";
		tbAddress  <="101001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111000101";
		tbAddress  <="101001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010001011";
		tbAddress  <="101001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100100011";
		tbAddress  <="101010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001010011";
		tbAddress  <="101010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010000011";
		tbAddress  <="101010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110000000";
		tbAddress  <="101010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111011111";
		tbAddress  <="101010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110010110";
		tbAddress  <="101010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001101001";
		tbAddress  <="101010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111001110";
		tbAddress  <="101010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010111011";
		tbAddress  <="101011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110000110";
		tbAddress  <="101011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110111100";
		tbAddress  <="101011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110101000";
		tbAddress  <="101011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010011110";
		tbAddress  <="101011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010110010";
		tbAddress  <="101011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000101110";
		tbAddress  <="101011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110001100";
		tbAddress  <="101011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100110110110";
		tbAddress  <="101100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011111011";
		tbAddress  <="101100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010101000";
		tbAddress  <="101100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100010001";
		tbAddress  <="101100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010101000";
		tbAddress  <="101100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111111100";
		tbAddress  <="101100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101101011";
		tbAddress  <="101100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100110110";
		tbAddress  <="101100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101100010";
		tbAddress  <="101101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011001001";
		tbAddress  <="101101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001110010";
		tbAddress  <="101101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101001101";
		tbAddress  <="101101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011100101";
		tbAddress  <="101101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000011110";
		tbAddress  <="101101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110111010";
		tbAddress  <="101101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000100000";
		tbAddress  <="101101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001011100";
		tbAddress  <="101110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110110110";
		tbAddress  <="101110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001100010";
		tbAddress  <="101110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000000101";
		tbAddress  <="101110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010111001";
		tbAddress  <="101110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001000000";
		tbAddress  <="101110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110100000";
		tbAddress  <="101110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110010011";
		tbAddress  <="101110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010011101";
		tbAddress  <="101111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111111";
		tbAddress  <="101111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000001010";
		tbAddress  <="101111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000110010";
		tbAddress  <="101111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010101011";
		tbAddress  <="101111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100111100";
		tbAddress  <="101111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001100000110";
		tbAddress  <="101111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111010111";
		tbAddress  <="101111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011111001";
		tbAddress  <="110000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111011001";
		tbAddress  <="110000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101001100";
		tbAddress  <="110000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110010011";
		tbAddress  <="110000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000011110";
		tbAddress  <="110000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011111110";
		tbAddress  <="110000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010001001";
		tbAddress  <="110000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110011010";
		tbAddress  <="110000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011001110";
		tbAddress  <="110001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011100001001";
		tbAddress  <="110001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000100110";
		tbAddress  <="110001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010101000";
		tbAddress  <="110001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001101111";
		tbAddress  <="110001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100000011";
		tbAddress  <="110001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011011101";
		tbAddress  <="110001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110011001100";
		tbAddress  <="110001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101100010";
		tbAddress  <="110010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110010110000";
		tbAddress  <="110010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001100001";
		tbAddress  <="110010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111000100";
		tbAddress  <="110010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110110101";
		tbAddress  <="110010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001001101";
		tbAddress  <="110010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001010010";
		tbAddress  <="110010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111001001";
		tbAddress  <="110010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111110111";
		tbAddress  <="110011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111010101";
		tbAddress  <="110011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100110000";
		tbAddress  <="110011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011010000";
		tbAddress  <="110011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010100001110";
		tbAddress  <="110011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100101111";
		tbAddress  <="110011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110110111";
		tbAddress  <="110011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110010";
		tbAddress  <="110011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010110110";
		tbAddress  <="110100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100110";
		tbAddress  <="110100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111101000";
		tbAddress  <="110100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000000010";
		tbAddress  <="110100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101001100";
		tbAddress  <="110100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101111111010";
		tbAddress  <="110100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110100110";
		tbAddress  <="110100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110110110";
		tbAddress  <="110100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111100011";
		tbAddress  <="110101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100111011";
		tbAddress  <="110101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101001111";
		tbAddress  <="110101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011101001";
		tbAddress  <="110101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011110010";
		tbAddress  <="110101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010000111";
		tbAddress  <="110101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010111110";
		tbAddress  <="110101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010110110";
		tbAddress  <="110101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100001111";
		tbAddress  <="110110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010100111";
		tbAddress  <="110110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000001101010";
		tbAddress  <="110110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101001001001";
		tbAddress  <="110110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011100011";
		tbAddress  <="110110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000110010";
		tbAddress  <="110110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110010010";
		tbAddress  <="110110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010111100";
		tbAddress  <="110110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101010011";
		tbAddress  <="110111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011001100";
		tbAddress  <="110111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010001011001";
		tbAddress  <="110111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110100000";
		tbAddress  <="110111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001101011";
		tbAddress  <="110111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101111100";
		tbAddress  <="110111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010111101";
		tbAddress  <="110111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101101101110";
		tbAddress  <="110111111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010101000";
		tbAddress  <="111000000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010100000";
		tbAddress  <="111000001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111010";
		tbAddress  <="111000010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001110011100";
		tbAddress  <="111000011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011011110";
		tbAddress  <="111000100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101010000101";
		tbAddress  <="111000101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010111110";
		tbAddress  <="111000110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100100100";
		tbAddress  <="111000111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001000011";
		tbAddress  <="111001000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110011101";
		tbAddress  <="111001001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111110000";
		tbAddress  <="111001010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010000011";
		tbAddress  <="111001011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000110100";
		tbAddress  <="111001100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000010111";
		tbAddress  <="111001101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011001110101";
		tbAddress  <="111001110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101011100111";
		tbAddress  <="111001111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000111111100";
		tbAddress  <="111010000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101001110";
		tbAddress  <="111010001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000111001";
		tbAddress  <="111010010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010001000";
		tbAddress  <="111010011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100101010110";
		tbAddress  <="111010100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000111011";
		tbAddress  <="111010101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110100010";
		tbAddress  <="111010110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010111100000";
		tbAddress  <="111010111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000000101";
		tbAddress  <="111011000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011011111";
		tbAddress  <="111011001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000000011010";
		tbAddress  <="111011010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100011111111";
		tbAddress  <="111011011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101001001";
		tbAddress  <="111011100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011101010";
		tbAddress  <="111011101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100010000101";
		tbAddress  <="111011110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110000001110";
		tbAddress  <="111011111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100110111";
		tbAddress  <="111100000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111000100";
		tbAddress  <="111100001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000010111011";
		tbAddress  <="111100010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="110001001101";
		tbAddress  <="111100011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011110000111";
		tbAddress  <="111100100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001011101100";
		tbAddress  <="111100101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000100001110";
		tbAddress  <="111100110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001101010110";
		tbAddress  <="111100111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100011001";
		tbAddress  <="111101000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101110011110";
		tbAddress  <="111101001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101000110000";
		tbAddress  <="111101010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010000100101";
		tbAddress  <="111101011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010110101001";
		tbAddress  <="111101100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101111111";
		tbAddress  <="111101101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100010001";
		tbAddress  <="111101110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011111010111";
		tbAddress  <="111101111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000101011000";
		tbAddress  <="111110000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100111110111";
		tbAddress  <="111110001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100100111110";
		tbAddress  <="111110010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001001110100";
		tbAddress  <="111110011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010011011100";
		tbAddress  <="111110100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011010000111";
		tbAddress  <="111110101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100111010";
		tbAddress  <="111110110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="101100001101";
		tbAddress  <="111110111";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000110001000";
		tbAddress  <="111111000";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010101000101";
		tbAddress  <="111111001";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="010010111110";
		tbAddress  <="111111010";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011000110101";
		tbAddress  <="111111011";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="011011111111";
		tbAddress  <="111111100";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="000011100000";
		tbAddress  <="111111101";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="100000110000";
		tbAddress  <="111111110";
		tbWE  <='1';
		wait for 10 ns;
		tbData_In  <="001010010010";
		tbAddress  <="111111111";
		tbWE  <='1';
		wait for 10 ns;
								
		tbWE  <='0';
		tbmode <= "01";
		tben<='1';
		
		wait for 10 ns;	
		
		tben<='0';
		
		wait for 30010 ns;	
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
		
	
END PROCESS;
	
  			
END test;
