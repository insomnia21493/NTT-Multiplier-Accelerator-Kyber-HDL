LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL; 
LIBRARY std;
USE std.standard.all;
LIBRARY work;
USE work.ALL;


ENTITY ntt IS

	PORT(
	
	clk         	:   IN  	std_logic;
	nrst        	:   IN  	std_logic;
	en	        	:   IN  	std_logic;
	mode	        :	IN		std_logic_vector(1 downto 0);
	
	WE				:	IN		std_logic;
	Address			:	IN		std_logic_vector(8 downto 0);
	Data_In			:	IN		std_logic_vector(11 downto 0);  
	Data_Out		:	OUT		std_logic_vector(11 downto 0);
	
	busy        	:   OUT 	std_logic;
	done        	:   OUT 	std_logic
	
	);


END ntt;




ARCHITECTURE behaviour OF ntt IS

--	attribute dont_touch : string;
--    attribute dont_touch of behaviour : architecture is "yes";

	 COMPONENT bf IS
					PORT(
				
				clk         :   IN 	std_logic;
				nrst        :   IN 	std_logic;
				
				bfmod		: 	IN  std_logic_vector(1 DOWNTO 0);
				
				rjin		: 	IN  std_logic_vector(11 DOWNTO 0);
				rjplin		: 	IN  std_logic_vector(11 DOWNTO 0);
				zeta 		: 	IN 	std_logic_vector(11 DOWNTO 0);
				
				rjout		: 	OUT std_logic_vector(11 DOWNTO 0);
				rjplout		: 	OUT std_logic_vector(11 DOWNTO 0)
				
				);

	 END COMPONENT;	
	 
	 

	 COMPONENT true_dpram_io IS
					PORT(
				
							clk			:	in		std_logic;
							we_a		:	in		std_logic;
							we_b		:	in		std_logic;
							data_a		:	in		std_logic_vector(11 downto 0);
							data_b		:	in		std_logic_vector(11 downto 0);
							addr_a		:	in		std_logic_vector(8 downto 0);
							addr_b		:	in		std_logic_vector(8 downto 0);
							q_a			:	out		std_logic_vector(11 downto 0);
							q_b			:	out		std_logic_vector(11 downto 0)
				
						);

	 END COMPONENT;	
	 
	 
	 COMPONENT true_dpram_temp1 IS
					PORT(
				
							clk			:	in		std_logic;
							we_a		:	in		std_logic;
							we_b		:	in		std_logic;
							data_a		:	in		std_logic_vector(11 downto 0);
							data_b		:	in		std_logic_vector(11 downto 0);
							addr_a		:	in		std_logic_vector(7 downto 0);
							addr_b		:	in		std_logic_vector(7 downto 0);
							q_a			:	out		std_logic_vector(11 downto 0);
							q_b			:	out		std_logic_vector(11 downto 0)
				
						);

	 END COMPONENT;	
	 
	 
	 COMPONENT true_dpram_temp2 IS
					PORT(
				
							clk			:	in		std_logic;
							we_a		:	in		std_logic;
							we_b		:	in		std_logic;
							data_a		:	in		std_logic_vector(11 downto 0);
							data_b		:	in		std_logic_vector(11 downto 0);
							addr_a		:	in		std_logic_vector(7 downto 0);
							addr_b		:	in		std_logic_vector(7 downto 0);
							q_a			:	out		std_logic_vector(11 downto 0);
							q_b			:	out		std_logic_vector(11 downto 0)
				
						);

	 END COMPONENT;	
	 
	 
	 COMPONENT ROM IS
					PORT(
				
							clk   : in std_logic;
							addr  : in std_logic_vector(7 downto 0);
							dout  : out std_logic_vector(11 downto 0)
							
							
						);

	 END COMPONENT;	
	 
	 
	TYPE state IS (idle , tontt, toinvntt , topwm );
	SIGNAL cur_st : state ;
	SIGNAL nxt_st : state;

	SIGNAL cntr		: std_logic_vector(11 downto 0);
	SIGNAL cntr1		: std_logic_vector(11 downto 0);
	
	SIGNAL iowea	: std_logic;
	SIGNAL ioweb	: std_logic;
	SIGNAL t1wea	: std_logic;
	SIGNAL t1web	: std_logic;
	SIGNAL t2wea	: std_logic;
	SIGNAL t2web	: std_logic;
	
	SIGNAL iodina	: std_logic_vector(11 downto 0);
	SIGNAL iodinb	: std_logic_vector(11 downto 0);
	SIGNAL iodouta	: std_logic_vector(11 downto 0);
	SIGNAL iodoutb	: std_logic_vector(11 downto 0);
	SIGNAL ioadda	: std_logic_vector(8 downto 0);
	SIGNAL ioaddb	: std_logic_vector(8 downto 0);
	SIGNAL t1dina	: std_logic_vector(11 downto 0);
	SIGNAL t1dinb	: std_logic_vector(11 downto 0);
	SIGNAL t1douta	: std_logic_vector(11 downto 0);
	SIGNAL t1doutb	: std_logic_vector(11 downto 0);
	SIGNAL t1adda	: std_logic_vector(7 downto 0);
	SIGNAL t1addb	: std_logic_vector(7 downto 0);
	SIGNAL t2dina	: std_logic_vector(11 downto 0);
	SIGNAL t2dinb	: std_logic_vector(11 downto 0);
	SIGNAL t2douta	: std_logic_vector(11 downto 0);
	SIGNAL t2doutb	: std_logic_vector(11 downto 0);
	SIGNAL t2adda	: std_logic_vector(7 downto 0);
	SIGNAL t2addb	: std_logic_vector(7 downto 0);
	
	SIGNAL zetain			    : unsigned(7 downto 0);
	SIGNAL zetaout			    : std_logic_vector(11 downto 0);
	SIGNAL bfmod		: std_logic_vector(1 DOWNTO 0);
	SIGNAL bfrjin		: std_logic_vector(11 DOWNTO 0);
	SIGNAL bfrjplin		: std_logic_vector(11 DOWNTO 0);
	SIGNAL bfzeta 		: std_logic_vector(11 DOWNTO 0);
	SIGNAL bfrjout		: std_logic_vector(11 DOWNTO 0);
	SIGNAL bfrjplout	: std_logic_vector(11 DOWNTO 0);
	
	SIGNAL wirebfrjout		: std_logic_vector(11 DOWNTO 0);
	SIGNAL wirebfrjplout	: std_logic_vector(11 DOWNTO 0);
	
	SIGNAL pdone	: std_logic;
	
	--attribute keep_hierarchy : string;
	--attribute keep_hierarchy of behaviour : ARCHITECTURE is "yes";
	
	attribute keep : string;
	
	attribute keep of iowea	 : signal is "true";
	attribute keep of ioweb	 : signal is "true";
	attribute keep of t1wea	 : signal is "true";
	attribute keep of t1web	 : signal is "true";
	attribute keep of t2wea	 : signal is "true";
	attribute keep of t2web	 : signal is "true";
	
	
	
	attribute keep of iodina	 : signal is "true";
	attribute keep of iodinb	 : signal is "true";
	--attribute keep of iodouta	 : signal is "true";
	--attribute keep of iodoutb	 : signal is "true";
	attribute keep of ioadda	 : signal is "true";
	attribute keep of ioaddb	 : signal is "true";
	attribute keep of t1dina	 : signal is "true";
	attribute keep of t1dinb	 : signal is "true";
	--attribute keep of t1douta	 : signal is "true";
	--attribute keep of t1doutb	 : signal is "true";
	attribute keep of t1adda	 : signal is "true";
	attribute keep of t1addb	 : signal is "true";
	attribute keep of t2dina	 : signal is "true";
	attribute keep of t2dinb	 : signal is "true";
	--attribute keep of t2douta	 : signal is "true";
	--attribute keep of t2doutb	 : signal is "true";
	attribute keep of t2adda	 : signal is "true";
	attribute keep of t2addb	 : signal is "true";
	
	attribute keep of wirebfrjout		 : signal is "true";
	attribute keep of wirebfrjplout	 : signal is "true";
	--
	--attribute dont_touch of cntr	 : signal is "true";
	--
	--
	--
	--attribute dont_touch of zetain		 : signal is "true";

	
	
	
	
	
	
	
	
	--attribute dont_touch of true_dpram_io : component is "yes";
	--attribute dont_touch of true_dpram_temp1 : component is "yes";
	--attribute dont_touch of true_dpram_temp2 : component is "yes";
	--attribute dont_touch of bf : component is "yes";
	
	
	
	
	
	
	
	
	
BEGIN


	bfc  :  bf PORT MAP(clk => clk , nrst => nrst ,  bfmod => bfmod , rjin => bfrjin  , rjplin => bfrjplin , zeta => bfzeta , rjout => wirebfrjout   , rjplout => wirebfrjplout   );

	ioram   :  true_dpram_io PORT MAP( clk => clk   , we_a =>  iowea  , we_b => ioweb , data_a => iodina   , data_b	=> iodinb   ,  addr_a	=>  ioadda , addr_b =>  ioaddb , q_a => iodouta , q_b =>  iodoutb  );
	temp1ram  :  true_dpram_temp1 PORT MAP( clk => clk  , we_a =>  t1wea  , we_b => t1web , data_a => t1dina   , data_b	=> t1dinb   ,  addr_a	=>  t1adda , addr_b =>  t1addb , q_a => t1douta , q_b =>  t1doutb  );
	temp2ram  :  true_dpram_temp2 PORT MAP( clk => clk  , we_a =>  t2wea  , we_b => t2web , data_a => t2dina   , data_b	=> t2dinb   ,  addr_a	=>  t2adda , addr_b =>  t2addb , q_a => t2douta , q_b =>  t2doutb  );
	
	zetarom: ROM PORT MAP( clk => clk , addr => std_logic_vector(zetain) , dout => zetaout);
	
		
	  bfzeta <= zetaout;



	

	
PROCESS(clk)
  BEGIN
  


  
  IF  clk'EVENT AND clk = '1' THEN
			
		IF nrst = '0' THEN

			cur_st<=idle;
			
			cntr <= "000000000000";
			
			
				iowea	<= '0';
				ioweb	<= '0';  
				t1wea	<= '0';  
				t1web	<= '0';  
				t2wea	<= '0';  
				t2web	<= '0';  
				pdone	<= '0';  
						
			--
				
				
				
				iodina		<= ( others => '0');
				iodinb	    <= ( others => '0');
				--iodouta	    <= ( others => '0');
				--iodoutb	    <= ( others => '0');
				ioadda	    <= ( others => '0');
				ioaddb	    <= ( others => '0');
				t1dina	    <= ( others => '0');
				t1dinb	    <= ( others => '0');
				--t1douta	    <= ( others => '0');
				--t1doutb	    <= ( others => '0');
				t1adda	    <= ( others => '0');
				t1addb	    <= ( others => '0');
				t2dina	    <= ( others => '0');
				t2dinb	    <= ( others => '0');
				--t2douta	    <= ( others => '0');
				--t2doutb	    <= ( others => '0');
				t2adda	    <= ( others => '0');
				t2addb	    <= ( others => '0');
				zetain	    <= ( others => '0');
				--zetaout	    <= ( others => '0');
				bfmod	    <= ( others => '0');
				bfrjin	    <= ( others => '0');
				bfrjplin	<= ( others => '0');
				--
				bfrjout	    <= ( others => '0');
				bfrjplout   <= ( others => '0');		

		ELSIF nrst='1' THEN
			
			cur_st <= nxt_st;
			
			pdone	<='0';
			
			iowea	<= '0';
			ioweb	<= '0';  
			t1wea	<= '0';  
			t1web	<= '0';  
			t2wea	<= '0';  
			t2web	<= '0';  
			
				cntr1 <= cntr;
	
	
	       bfrjout		<= wirebfrjout	;
            bfrjplout   <= wirebfrjplout;
		
			IF cur_st = idle THEN
				
				cntr <= "000000000000";
				cntr1 <= "000000000000";
				
				iowea <= WE;
				ioadda <= Address;
				iodina <= Data_In;
				Data_Out <= iodouta;
				

			
			ELSIF cur_st = tontt THEN
				
				IF cntr = "000000000000" THEN
					
					ioadda <= "000000000";
					ioaddb <= "010000000";
					
					bfmod <= "00";
					
					zetain <= "00000001";
					
					cntr <= "000000000001";
				
				ELSIF cntr = "000000000001" THEN
				
					ioadda <= "000000001";
					ioaddb <= "010000001";
					
					
					cntr <= "000000000010";
					
				ELSIF cntr = "000000000010" THEN
					
					ioadda <= "000000010";
					ioaddb <= "010000010";
					
					bfrjin 	 <= iodouta;
					bfrjplin <= iodoutb;
					
					
					
					cntr <= "000000000011";
				
				ELSIF cntr = "000000000011" THEN
				
					ioadda <= "000000011";
					ioaddb <= "010000011";
					
					bfrjin 	 <= iodouta;
					bfrjplin <= iodoutb;
					
					cntr <= "000000000100";
					
				ELSIF cntr = "000000000100" THEN
					
					ioadda <= "000000100";
					ioaddb <= "010000100";
					
					bfrjin 	 <= iodouta;
					bfrjplin <= iodoutb;
				
					cntr <= "000000000101";
				
				ELSIF cntr = "000000000101" THEN
					
					ioadda <= "000000101";
					ioaddb <= "010000101";
				
					bfrjin 	 <= iodouta;
					bfrjplin <= iodoutb;
					
					cntr <= "000000000110";
				
				ELSIF cntr = "000000000110" THEN
				
					ioadda <= "000000110";
					ioaddb <= "010000110";
					
					bfrjin 	 <= iodouta;
					bfrjplin <= iodoutb;
					
					
					
					
					cntr <= "000000000111";
				elsif cntr ="000000000111" THEN
				      ioadda <= "000000111";
				      ioaddb <= "010000111";
				
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				      cntr <= "000000001000";
				elsif cntr ="000000001000" THEN
				      ioadda <= "000001000";
				      ioaddb <= "010001000";
				
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				      cntr <= "000000001001";
				elsif cntr ="000000001001" THEN
				      ioadda <= "000001001";
				      ioaddb <= "010001001";
				
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
					  	  					  
				      cntr <= "000000001010";
				elsif cntr ="000000001010" THEN
				      ioadda <= "000001010";
				      ioaddb <= "010001010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000001011";
				elsif cntr ="000000001011" THEN
				      ioadda <= "000001011";
				      ioaddb <= "010001011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000001100";
				elsif cntr ="000000001100" THEN
				      ioadda <= "000001100";
				      ioaddb <= "010001100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000001101";
				elsif cntr ="000000001101" THEN
				      ioadda <= "000001101";
				      ioaddb <= "010001101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000001110";
				elsif cntr ="000000001110" THEN
				      ioadda <= "000001110";
				      ioaddb <= "010001110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000001111";
				elsif cntr ="000000001111" THEN
				      ioadda <= "000001111";
				      ioaddb <= "010001111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010000";
				elsif cntr ="000000010000" THEN
				      ioadda <= "000010000";
				      ioaddb <= "010010000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010001";
				elsif cntr ="000000010001" THEN
				      ioadda <= "000010001";
				      ioaddb <= "010010001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010010";
				elsif cntr ="000000010010" THEN
				      ioadda <= "000010010";
				      ioaddb <= "010010010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010011";
				elsif cntr ="000000010011" THEN
				      ioadda <= "000010011";
				      ioaddb <= "010010011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010100";
				elsif cntr ="000000010100" THEN
				      ioadda <= "000010100";
				      ioaddb <= "010010100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010101";
				elsif cntr ="000000010101" THEN
				      ioadda <= "000010101";
				      ioaddb <= "010010101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010110";
				elsif cntr ="000000010110" THEN
				      ioadda <= "000010110";
				      ioaddb <= "010010110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000010111";
				elsif cntr ="000000010111" THEN
				      ioadda <= "000010111";
				      ioaddb <= "010010111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011000";
				elsif cntr ="000000011000" THEN
				      ioadda <= "000011000";
				      ioaddb <= "010011000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011001";
				elsif cntr ="000000011001" THEN
				      ioadda <= "000011001";
				      ioaddb <= "010011001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011010";
				elsif cntr ="000000011010" THEN
				      ioadda <= "000011010";
				      ioaddb <= "010011010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011011";
				elsif cntr ="000000011011" THEN
				      ioadda <= "000011011";
				      ioaddb <= "010011011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011100";
				elsif cntr ="000000011100" THEN
				      ioadda <= "000011100";
				      ioaddb <= "010011100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011101";
				elsif cntr ="000000011101" THEN
				      ioadda <= "000011101";
				      ioaddb <= "010011101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011110";
				elsif cntr ="000000011110" THEN
				      ioadda <= "000011110";
				      ioaddb <= "010011110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000011111";
				elsif cntr ="000000011111" THEN
				      ioadda <= "000011111";
				      ioaddb <= "010011111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100000";
				elsif cntr ="000000100000" THEN
				      ioadda <= "000100000";
				      ioaddb <= "010100000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100001";
				elsif cntr ="000000100001" THEN
				      ioadda <= "000100001";
				      ioaddb <= "010100001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100010";
				elsif cntr ="000000100010" THEN
				      ioadda <= "000100010";
				      ioaddb <= "010100010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100011";
				elsif cntr ="000000100011" THEN
				      ioadda <= "000100011";
				      ioaddb <= "010100011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100100";
				elsif cntr ="000000100100" THEN
				      ioadda <= "000100100";
				      ioaddb <= "010100100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100101";
				elsif cntr ="000000100101" THEN
				      ioadda <= "000100101";
				      ioaddb <= "010100101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100110";
				elsif cntr ="000000100110" THEN
				      ioadda <= "000100110";
				      ioaddb <= "010100110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000100111";
				elsif cntr ="000000100111" THEN
				      ioadda <= "000100111";
				      ioaddb <= "010100111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101000";
				elsif cntr ="000000101000" THEN
				      ioadda <= "000101000";
				      ioaddb <= "010101000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101001";
				elsif cntr ="000000101001" THEN
				      ioadda <= "000101001";
				      ioaddb <= "010101001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101010";
				elsif cntr ="000000101010" THEN
				      ioadda <= "000101010";
				      ioaddb <= "010101010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101011";
				elsif cntr ="000000101011" THEN
				      ioadda <= "000101011";
				      ioaddb <= "010101011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101100";
				elsif cntr ="000000101100" THEN
				      ioadda <= "000101100";
				      ioaddb <= "010101100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101101";
				elsif cntr ="000000101101" THEN
				      ioadda <= "000101101";
				      ioaddb <= "010101101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101110";
				elsif cntr ="000000101110" THEN
				      ioadda <= "000101110";
				      ioaddb <= "010101110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000101111";
				elsif cntr ="000000101111" THEN
				      ioadda <= "000101111";
				      ioaddb <= "010101111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110000";
				elsif cntr ="000000110000" THEN
				      ioadda <= "000110000";
				      ioaddb <= "010110000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110001";
				elsif cntr ="000000110001" THEN
				      ioadda <= "000110001";
				      ioaddb <= "010110001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110010";
				elsif cntr ="000000110010" THEN
				      ioadda <= "000110010";
				      ioaddb <= "010110010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110011";
				elsif cntr ="000000110011" THEN
				      ioadda <= "000110011";
				      ioaddb <= "010110011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110100";
				elsif cntr ="000000110100" THEN
				      ioadda <= "000110100";
				      ioaddb <= "010110100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110101";
				elsif cntr ="000000110101" THEN
				      ioadda <= "000110101";
				      ioaddb <= "010110101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110110";
				elsif cntr ="000000110110" THEN
				      ioadda <= "000110110";
				      ioaddb <= "010110110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000110111";
				elsif cntr ="000000110111" THEN
				      ioadda <= "000110111";
				      ioaddb <= "010110111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111000";
				elsif cntr ="000000111000" THEN
				      ioadda <= "000111000";
				      ioaddb <= "010111000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111001";
				elsif cntr ="000000111001" THEN
				      ioadda <= "000111001";
				      ioaddb <= "010111001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111010";
				elsif cntr ="000000111010" THEN
				      ioadda <= "000111010";
				      ioaddb <= "010111010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111011";
				elsif cntr ="000000111011" THEN
				      ioadda <= "000111011";
				      ioaddb <= "010111011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111100";
				elsif cntr ="000000111100" THEN
				      ioadda <= "000111100";
				      ioaddb <= "010111100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111101";
				elsif cntr ="000000111101" THEN
				      ioadda <= "000111101";
				      ioaddb <= "010111101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111110";
				elsif cntr ="000000111110" THEN
				      ioadda <= "000111110";
				      ioaddb <= "010111110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000000111111";
				elsif cntr ="000000111111" THEN
				      ioadda <= "000111111";
				      ioaddb <= "010111111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000000";
				elsif cntr ="000001000000" THEN
				      ioadda <= "001000000";
				      ioaddb <= "011000000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000001";
				elsif cntr ="000001000001" THEN
				      ioadda <= "001000001";
				      ioaddb <= "011000001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000010";
				elsif cntr ="000001000010" THEN
				      ioadda <= "001000010";
				      ioaddb <= "011000010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000011";
				elsif cntr ="000001000011" THEN
				      ioadda <= "001000011";
				      ioaddb <= "011000011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000100";
				elsif cntr ="000001000100" THEN
				      ioadda <= "001000100";
				      ioaddb <= "011000100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000101";
				elsif cntr ="000001000101" THEN
				      ioadda <= "001000101";
				      ioaddb <= "011000101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000110";
				elsif cntr ="000001000110" THEN
				      ioadda <= "001000110";
				      ioaddb <= "011000110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001000111";
				elsif cntr ="000001000111" THEN
				      ioadda <= "001000111";
				      ioaddb <= "011000111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001000";
				elsif cntr ="000001001000" THEN
				      ioadda <= "001001000";
				      ioaddb <= "011001000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001001";
				elsif cntr ="000001001001" THEN
				      ioadda <= "001001001";
				      ioaddb <= "011001001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001010";
				elsif cntr ="000001001010" THEN
				      ioadda <= "001001010";
				      ioaddb <= "011001010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001011";
				elsif cntr ="000001001011" THEN
				      ioadda <= "001001011";
				      ioaddb <= "011001011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001100";
				elsif cntr ="000001001100" THEN
				      ioadda <= "001001100";
				      ioaddb <= "011001100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001101";
				elsif cntr ="000001001101" THEN
				      ioadda <= "001001101";
				      ioaddb <= "011001101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001110";
				elsif cntr ="000001001110" THEN
				      ioadda <= "001001110";
				      ioaddb <= "011001110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001001111";
				elsif cntr ="000001001111" THEN
				      ioadda <= "001001111";
				      ioaddb <= "011001111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010000";
				elsif cntr ="000001010000" THEN
				      ioadda <= "001010000";
				      ioaddb <= "011010000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010001";
				elsif cntr ="000001010001" THEN
				      ioadda <= "001010001";
				      ioaddb <= "011010001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010010";
				elsif cntr ="000001010010" THEN
				      ioadda <= "001010010";
				      ioaddb <= "011010010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010011";
				elsif cntr ="000001010011" THEN
				      ioadda <= "001010011";
				      ioaddb <= "011010011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010100";
				elsif cntr ="000001010100" THEN
				      ioadda <= "001010100";
				      ioaddb <= "011010100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010101";
				elsif cntr ="000001010101" THEN
				      ioadda <= "001010101";
				      ioaddb <= "011010101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010110";
				elsif cntr ="000001010110" THEN
				      ioadda <= "001010110";
				      ioaddb <= "011010110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001010111";
				elsif cntr ="000001010111" THEN
				      ioadda <= "001010111";
				      ioaddb <= "011010111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011000";
				elsif cntr ="000001011000" THEN
				      ioadda <= "001011000";
				      ioaddb <= "011011000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011001";
				elsif cntr ="000001011001" THEN
				      ioadda <= "001011001";
				      ioaddb <= "011011001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011010";
				elsif cntr ="000001011010" THEN
				      ioadda <= "001011010";
				      ioaddb <= "011011010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011011";
				elsif cntr ="000001011011" THEN
				      ioadda <= "001011011";
				      ioaddb <= "011011011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011100";
				elsif cntr ="000001011100" THEN
				      ioadda <= "001011100";
				      ioaddb <= "011011100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011101";
				elsif cntr ="000001011101" THEN
				      ioadda <= "001011101";
				      ioaddb <= "011011101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011110";
				elsif cntr ="000001011110" THEN
				      ioadda <= "001011110";
				      ioaddb <= "011011110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001011111";
				elsif cntr ="000001011111" THEN
				      ioadda <= "001011111";
				      ioaddb <= "011011111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100000";
				elsif cntr ="000001100000" THEN
				      ioadda <= "001100000";
				      ioaddb <= "011100000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100001";
				elsif cntr ="000001100001" THEN
				      ioadda <= "001100001";
				      ioaddb <= "011100001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100010";
				elsif cntr ="000001100010" THEN
				      ioadda <= "001100010";
				      ioaddb <= "011100010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100011";
				elsif cntr ="000001100011" THEN
				      ioadda <= "001100011";
				      ioaddb <= "011100011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100100";
				elsif cntr ="000001100100" THEN
				      ioadda <= "001100100";
				      ioaddb <= "011100100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100101";
				elsif cntr ="000001100101" THEN
				      ioadda <= "001100101";
				      ioaddb <= "011100101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100110";
				elsif cntr ="000001100110" THEN
				      ioadda <= "001100110";
				      ioaddb <= "011100110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001100111";
				elsif cntr ="000001100111" THEN
				      ioadda <= "001100111";
				      ioaddb <= "011100111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101000";
				elsif cntr ="000001101000" THEN
				      ioadda <= "001101000";
				      ioaddb <= "011101000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101001";
				elsif cntr ="000001101001" THEN
				      ioadda <= "001101001";
				      ioaddb <= "011101001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101010";
				elsif cntr ="000001101010" THEN
				      ioadda <= "001101010";
				      ioaddb <= "011101010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101011";
				elsif cntr ="000001101011" THEN
				      ioadda <= "001101011";
				      ioaddb <= "011101011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101100";
				elsif cntr ="000001101100" THEN
				      ioadda <= "001101100";
				      ioaddb <= "011101100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101101";
				elsif cntr ="000001101101" THEN
				      ioadda <= "001101101";
				      ioaddb <= "011101101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101110";
				elsif cntr ="000001101110" THEN
				      ioadda <= "001101110";
				      ioaddb <= "011101110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001101111";
				elsif cntr ="000001101111" THEN
				      ioadda <= "001101111";
				      ioaddb <= "011101111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110000";
				elsif cntr ="000001110000" THEN
				      ioadda <= "001110000";
				      ioaddb <= "011110000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110001";
				elsif cntr ="000001110001" THEN
				      ioadda <= "001110001";
				      ioaddb <= "011110001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110010";
				elsif cntr ="000001110010" THEN
				      ioadda <= "001110010";
				      ioaddb <= "011110010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110011";
				elsif cntr ="000001110011" THEN
				      ioadda <= "001110011";
				      ioaddb <= "011110011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110100";
				elsif cntr ="000001110100" THEN
				      ioadda <= "001110100";
				      ioaddb <= "011110100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110101";
				elsif cntr ="000001110101" THEN
				      ioadda <= "001110101";
				      ioaddb <= "011110101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110110";
				elsif cntr ="000001110110" THEN
				      ioadda <= "001110110";
				      ioaddb <= "011110110";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001110111";
				elsif cntr ="000001110111" THEN
				      ioadda <= "001110111";
				      ioaddb <= "011110111";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111000";
				elsif cntr ="000001111000" THEN
				      ioadda <= "001111000";
				      ioaddb <= "011111000";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111001";
				elsif cntr ="000001111001" THEN
				      ioadda <= "001111001";
				      ioaddb <= "011111001";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111010";
				elsif cntr ="000001111010" THEN
				      ioadda <= "001111010";
				      ioaddb <= "011111010";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111011";
				elsif cntr ="000001111011" THEN
				      ioadda <= "001111011";
				      ioaddb <= "011111011";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111100";
				elsif cntr ="000001111100" THEN
				      ioadda <= "001111100";
				      ioaddb <= "011111100";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111101";
				elsif cntr ="000001111101" THEN
				      ioadda <= "001111101";
				      ioaddb <= "011111101";
				      
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111110";
				elsif cntr ="000001111110" THEN
				      ioadda <= "001111110";
				      ioaddb <= "011111110";
				      
					  
					 
					  
					  
					  
					  
					  
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000001111111";
				elsif cntr ="000001111111" THEN
				      ioadda <= "001111111";
				      ioaddb <= "011111111";
				      
					  
					  
					  
					  
					  
					  
					  
					  
				      bfrjin     <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      cntr <= "000010000000";
				elsif cntr ="000010000000" THEN
				      
					  t1addb <= "00000000";
					  t2addb <= "01000000";
					  
					  
					  
					  bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
					  
				      
				      
					  cntr <= "000010000001";
				elsif cntr ="000010000001" THEN
					  
					  t1addb <= "00000001";
					  t2addb <= "01000001";
					  
					  zetain   <="00000010";
					  
					  bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
					  
					  
					  
					  cntr <= "000010000010";
				elsif cntr ="000010000010" THEN
					  
					  t1addb <= "00000010";
				      t2addb <= "01000010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;

					  
					  
					  
					  
					  cntr <= "000010000011";
				elsif cntr ="000010000011" THEN
					  
					       t1addb <= "00000011";
      t2addb <= "01000011";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb; 
					  
					  
					  
					  
					  cntr <= "000010000100";
				elsif cntr ="000010000100" THEN
					  
					  
					  t1addb <= "00000100";
      t2addb <= "01000100";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb;
					  
					  
					  
					  cntr <= "000010000101";
				elsif cntr ="000010000101" THEN
					  
					   t1addb <= "00000101";
      t2addb <= "01000101";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb;
					  
					  
					  
					  
					  cntr <= "000010000110";
				elsif cntr ="000010000110" THEN
					  
					  t1addb <= "00000110";
      t2addb <= "01000110";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb;

					  
					  
					  
					  
					  cntr <= "000010000111";
				elsif cntr ="000010000111" THEN
					  
					  t1addb <= "00000111";
      t2addb <= "01000111";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb;

					  
					  
					  
					  
					  cntr <= "000010001000";
				elsif cntr ="000010001000" THEN
					  
					  t1addb <= "00001000";
      t2addb <= "01001000";
      bfrjin     <= t1doutb;
      bfrjplin <= t2doutb;



					  
					  
					  
					  
					  cntr <= "000010001001";
				elsif cntr ="000010001001" THEN
				      t1addb <= "00001001";
				      t2addb <= "01001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
					  
				      
				      
				      
				      cntr <= "000010001010";
				elsif cntr ="000010001010" THEN
				      t1addb <= "00001010";  
				      t2addb <= "01001010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010001011";  
				elsif cntr ="000010001011" THEN
				      t1addb <= "00001011";
				      t2addb <= "01001011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010001100";
				elsif cntr ="000010001100" THEN
				      t1addb <= "00001100";
				      t2addb <= "01001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010001101";
				elsif cntr ="000010001101" THEN
				      t1addb <= "00001101";
				      t2addb <= "01001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010001110";
				elsif cntr ="000010001110" THEN
				      t1addb <= "00001110";
				      t2addb <= "01001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010001111";
				elsif cntr ="000010001111" THEN
				      t1addb <= "00001111";
				      t2addb <= "01001111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
				      
				      cntr <= "000010010000";
				elsif cntr ="000010010000" THEN
				      t1addb <= "00010000";  
				      t2addb <= "01010000";  
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010001";
				elsif cntr ="000010010001" THEN
				      t1addb <= "00010001";
				      t2addb <= "01010001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010010";
				elsif cntr ="000010010010" THEN
				      t1addb <= "00010010";
				      t2addb <= "01010010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010011";  
				elsif cntr ="000010010011" THEN
				      t1addb <= "00010011";
				      t2addb <= "01010011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010100";
				elsif cntr ="000010010100" THEN
				      t1addb <= "00010100";
				      t2addb <= "01010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010101";
				elsif cntr ="000010010101" THEN
				      t1addb <= "00010101";
				      t2addb <= "01010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010110";
				elsif cntr ="000010010110" THEN
				      t1addb <= "00010110";
				      t2addb <= "01010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010010111";
				elsif cntr ="000010010111" THEN
				      t1addb <= "00010111";
				      t2addb <= "01010111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
				      
				      cntr <= "000010011000";
				elsif cntr ="000010011000" THEN
				      t1addb <= "00011000";  
				      t2addb <= "01011000";  
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011001";  
				elsif cntr ="000010011001" THEN  
				      t1addb <= "00011001";
				      t2addb <= "01011001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011010";
				elsif cntr ="000010011010" THEN
				      t1addb <= "00011010";  
				      t2addb <= "01011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011011";
				elsif cntr ="000010011011" THEN
				      t1addb <= "00011011";
				      t2addb <= "01011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011100";
				elsif cntr ="000010011100" THEN
				      t1addb <= "00011100";
				      t2addb <= "01011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011101";
				elsif cntr ="000010011101" THEN
				      t1addb <= "00011101";
				      t2addb <= "01011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011110";
				elsif cntr ="000010011110" THEN
				      t1addb <= "00011110";
				      t2addb <= "01011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010011111";
				elsif cntr ="000010011111" THEN
				      t1addb <= "00011111";
				      t2addb <= "01011111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
				      
				      cntr <= "000010100000";
				elsif cntr ="000010100000" THEN
				      t1addb <= "00100000";  
				      t2addb <= "01100000";  
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100001";  
				elsif cntr ="000010100001" THEN  
				      t1addb <= "00100001";
				      t2addb <= "01100001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100010";
				elsif cntr ="000010100010" THEN
				      t1addb <= "00100010";  
				      t2addb <= "01100010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100011";  
				elsif cntr ="000010100011" THEN
				      t1addb <= "00100011";
				      t2addb <= "01100011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100100";
				elsif cntr ="000010100100" THEN
				      t1addb <= "00100100";
				      t2addb <= "01100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100101";
				elsif cntr ="000010100101" THEN
				      t1addb <= "00100101";
				      t2addb <= "01100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100110";
				elsif cntr ="000010100110" THEN
				      t1addb <= "00100110";
				      t2addb <= "01100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010100111";
				elsif cntr ="000010100111" THEN
				      t1addb <= "00100111";
				      t2addb <= "01100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101000";
				elsif cntr ="000010101000" THEN
				      t1addb <= "00101000";  
				      t2addb <= "01101000";  
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101001";  
				elsif cntr ="000010101001" THEN  
				      t1addb <= "00101001";
				      t2addb <= "01101001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101010";
				elsif cntr ="000010101010" THEN
				      t1addb <= "00101010";  
				      t2addb <= "01101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101011";  
				elsif cntr ="000010101011" THEN
				      t1addb <= "00101011";
				      t2addb <= "01101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101100";
				elsif cntr ="000010101100" THEN
				      t1addb <= "00101100";
				      t2addb <= "01101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101101";
				elsif cntr ="000010101101" THEN
				      t1addb <= "00101101";
				      t2addb <= "01101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101110";
				elsif cntr ="000010101110" THEN
				      t1addb <= "00101110";
				      t2addb <= "01101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010101111";
				elsif cntr ="000010101111" THEN
				      t1addb <= "00101111";
				      t2addb <= "01101111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
				      
				      cntr <= "000010110000";
				elsif cntr ="000010110000" THEN
				      t1addb <= "00110000";
				      t2addb <= "01110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110001";  
				elsif cntr ="000010110001" THEN  
				      t1addb <= "00110001";
				      t2addb <= "01110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110010";
				elsif cntr ="000010110010" THEN
				      t1addb <= "00110010";  
				      t2addb <= "01110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110011";  
				elsif cntr ="000010110011" THEN
				      t1addb <= "00110011";
				      t2addb <= "01110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110100";
				elsif cntr ="000010110100" THEN
				      t1addb <= "00110100";
				      t2addb <= "01110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110101";
				elsif cntr ="000010110101" THEN
				      t1addb <= "00110101";
				      t2addb <= "01110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110110";
				elsif cntr ="000010110110" THEN
				      t1addb <= "00110110";
				      t2addb <= "01110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010110111";
				elsif cntr ="000010110111" THEN
				      t1addb <= "00110111";
				      t2addb <= "01110111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
				      
				      cntr <= "000010111000";
				elsif cntr ="000010111000" THEN
				      t1addb <= "00111000";  
				      t2addb <= "01111000";  
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111001";
				elsif cntr ="000010111001" THEN
				      t1addb <= "00111001";
				      t2addb <= "01111001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111010";
				elsif cntr ="000010111010" THEN
				      t1addb <= "00111010";
				      t2addb <= "01111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111011";  
				elsif cntr ="000010111011" THEN
				      t1addb <= "00111011";
				      t2addb <= "01111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111100";
				elsif cntr ="000010111100" THEN
				      t1addb <= "00111100";
				      t2addb <= "01111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111101";
				elsif cntr ="000010111101" THEN
				      t1addb <= "00111101";
				      t2addb <= "01111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111110";
				elsif cntr ="000010111110" THEN
				      t1addb <= "00111110";
				      t2addb <= "01111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000010111111";
				elsif cntr ="000010111111" THEN
				      t1addb <= "00111111";
				      t2addb <= "01111111";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb;  
				      
				      
				      
					  
				      cntr <= "000011000000";
				elsif cntr ="000011000000" THEN
				      t1addb <= "01000000";  
				      t2addb <= "00000000";  
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb; 
				      
				      
				      
				      
				      cntr <= "000011000001";  
				elsif cntr ="000011000001" THEN  
				      t1addb <= "01000001";
				      t2addb <= "00000001";
				      bfrjin     <= t1doutb;  
				      bfrjplin <= t2doutb; 
				      
				      
				      
					  zetain   <="00000011";
				      cntr <= "000011000010";
				elsif cntr ="000011000010" THEN
				      t1addb <= "01000010";  
				      t2addb <= "00000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
					  
					  
				      cntr <= "000011000011";
				elsif cntr ="000011000011" THEN
				      t1addb <= "01000011";
				      t2addb <= "00000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011000100";
				elsif cntr ="000011000100" THEN
				      t1addb <= "01000100";
				      t2addb <= "00000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011000101";
				elsif cntr ="000011000101" THEN
				      t1addb <= "01000101";
				      t2addb <= "00000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011000110";
				elsif cntr ="000011000110" THEN
				      t1addb <= "01000110";
				      t2addb <= "00000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011000111";
				elsif cntr ="000011000111" THEN
				      t1addb <= "01000111";
				      t2addb <= "00000111";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;  
				      
				      
				      
				      
				      cntr <= "000011001000";
				elsif cntr ="000011001000" THEN
				      t1addb <= "01001000";  
				      t2addb <= "00001000";  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001001";  
				elsif cntr ="000011001001" THEN  
				      t1addb <= "01001001";
				      t2addb <= "00001001";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001010";
				elsif cntr ="000011001010" THEN
				      t1addb <= "01001010";  
				      t2addb <= "00001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001011";  
				elsif cntr ="000011001011" THEN
				      t1addb <= "01001011";
				      t2addb <= "00001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001100";
				elsif cntr ="000011001100" THEN
				      t1addb <= "01001100";
				      t2addb <= "00001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001101";
				elsif cntr ="000011001101" THEN
				      t1addb <= "01001101";
				      t2addb <= "00001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001110";
				elsif cntr ="000011001110" THEN
				      t1addb <= "01001110";
				      t2addb <= "00001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011001111";
				elsif cntr ="000011001111" THEN
				      t1addb <= "01001111";
				      t2addb <= "00001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010000";
				elsif cntr ="000011010000" THEN
				      t1addb <= "01010000";  
				      t2addb <= "00010000";  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010001";  
				elsif cntr ="000011010001" THEN  
				      t1addb <= "01010001";
				      t2addb <= "00010001";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010010";
				elsif cntr ="000011010010" THEN
				      t1addb <= "01010010";  
				      t2addb <= "00010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010011";  
				elsif cntr ="000011010011" THEN
				      t1addb <= "01010011";
				      t2addb <= "00010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010100";
				elsif cntr ="000011010100" THEN
				      t1addb <= "01010100";
				      t2addb <= "00010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010101";
				elsif cntr ="000011010101" THEN
				      t1addb <= "01010101";
				      t2addb <= "00010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010110";
				elsif cntr ="000011010110" THEN
				      t1addb <= "01010110";
				      t2addb <= "00010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011010111";
				elsif cntr ="000011010111" THEN
				      t1addb <= "01010111";
				      t2addb <= "00010111";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;  
				      
				      
				      
				      
				      cntr <= "000011011000";
				elsif cntr ="000011011000" THEN
				      t1addb <= "01011000";
				      t2addb <= "00011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011001";  
				elsif cntr ="000011011001" THEN  
				      t1addb <= "01011001";
				      t2addb <= "00011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011010";
				elsif cntr ="000011011010" THEN
				      t1addb <= "01011010";  
				      t2addb <= "00011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011011";  
				elsif cntr ="000011011011" THEN
				      t1addb <= "01011011";
				      t2addb <= "00011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011100";
				elsif cntr ="000011011100" THEN
				      t1addb <= "01011100";
				      t2addb <= "00011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011101";
				elsif cntr ="000011011101" THEN
				      t1addb <= "01011101";
				      t2addb <= "00011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011110";
				elsif cntr ="000011011110" THEN
				      t1addb <= "01011110";
				      t2addb <= "00011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011011111";
				elsif cntr ="000011011111" THEN
				      t1addb <= "01011111";
				      t2addb <= "00011111";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;  
				      
				      
				      
				      
				      cntr <= "000011100000";
				elsif cntr ="000011100000" THEN
				      t1addb <= "01100000";  
				      t2addb <= "00100000";  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100001";
				elsif cntr ="000011100001" THEN
				      t1addb <= "01100001";
				      t2addb <= "00100001";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100010";
				elsif cntr ="000011100010" THEN
				      t1addb <= "01100010";
				      t2addb <= "00100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100011";  
				elsif cntr ="000011100011" THEN
				      t1addb <= "01100011";
				      t2addb <= "00100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100100";
				elsif cntr ="000011100100" THEN
				      t1addb <= "01100100";
				      t2addb <= "00100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100101";
				elsif cntr ="000011100101" THEN
				      t1addb <= "01100101";
				      t2addb <= "00100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100110";
				elsif cntr ="000011100110" THEN
				      t1addb <= "01100110";
				      t2addb <= "00100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011100111";
				elsif cntr ="000011100111" THEN
				      t1addb <= "01100111";
				      t2addb <= "00100111";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;  
				      
				      
				      
				      
				      cntr <= "000011101000";
				elsif cntr ="000011101000" THEN
				      t1addb <= "01101000";  
				      t2addb <= "00101000";  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101001";  
				elsif cntr ="000011101001" THEN  
				      t1addb <= "01101001";
				      t2addb <= "00101001";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;
				      
				      
				      
			          
				      cntr <= "000011101010";
				elsif cntr ="000011101010" THEN
				      t1addb <= "01101010";  
				      t2addb <= "00101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101011";  
				elsif cntr ="000011101011" THEN
				      t1addb <= "01101011";
				      t2addb <= "00101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101100";
				elsif cntr ="000011101100" THEN
				      t1addb <= "01101100";
				      t2addb <= "00101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101101";
				elsif cntr ="000011101101" THEN
				      t1addb <= "01101101";
				      t2addb <= "00101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101110";
				elsif cntr ="000011101110" THEN
				      t1addb <= "01101110";
				      t2addb <= "00101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011101111";
				elsif cntr ="000011101111" THEN
				      t1addb <= "01101111";
				      t2addb <= "00101111";
				      bfrjin     <= t2doutb;  
				      bfrjplin <= t1doutb;  
				      
				      
				      
				      
				      cntr <= "000011110000";
				elsif cntr ="000011110000" THEN
				      t1addb <= "01110000";
				      t2addb <= "00110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011110001";  
				elsif cntr ="000011110001" THEN  
				      t1addb <= "01110001";
				      t2addb <= "00110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011110010";
				elsif cntr ="000011110010" THEN
				      t1addb <= "01110010";  
				      t2addb <= "00110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000011110011";
				elsif cntr ="000011110011" THEN
				      t1addb <= "01110011";
				      t2addb <= "00110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011110100";
				elsif cntr ="000011110100" THEN
				      t1addb <= "01110100";	  
				      t2addb <= "00110100";	  
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011110101";	  
				elsif cntr ="000011110101" THEN	  
				      t1addb <= "01110101";
				      t2addb <= "00110101";
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011110110";	  
				elsif cntr ="000011110110" THEN	  
				      t1addb <= "01110110";	  
				      t2addb <= "00110110";	  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
					  
				      
					  
					  
				      cntr <= "000011110111";	  
				elsif cntr ="000011110111" THEN	  
				      t1addb <= "01110111";	  
				      t2addb <= "00110111";	  
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
				      
					  
				      
				      
				      cntr <= "000011111000";	  
				elsif cntr ="000011111000" THEN	  
				      t1addb <= "01111000";	  
				      t2addb <= "00111000";	  
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011111001";
				elsif cntr ="000011111001" THEN
				      t1addb <= "01111001";	  
				      t2addb <= "00111001";	  
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011111010";	  
				elsif cntr ="000011111010" THEN	  
				      t1addb <= "01111010";
				      t2addb <= "00111010";
				      bfrjin     <= t2doutb;	  
				      bfrjplin <= t1doutb;	  
					  
					  
					  
					  
				      cntr <= "000011111011";	  
				elsif cntr ="000011111011" THEN	  
				      t1addb <= "01111011";	  
				      t2addb <= "00111011";	  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
					  
					  
					  
					  
				      cntr <= "000011111100";	  
				elsif cntr ="000011111100" THEN	  
				      t1addb <= "01111100";	  
				      t2addb <= "00111100";	  
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
					  
                      
                      
                      
                      cntr <= "000011111101";
                elsif cntr ="000011111101" THEN
                      t1addb <= "01111101";
                      t2addb <= "00111101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "000011111110";
                elsif cntr ="000011111110" THEN
                      t1addb <= "01111110";
                      t2addb <= "00111110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      cntr <= "000011111111";
                elsif cntr ="000011111111" THEN
                      t1addb <= "01111111";
                      t2addb <= "00111111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      cntr <= "000100000000";
				elsif cntr ="000100000000" THEN
				      t1addb <= "10000000";
				      t2addb <= "10100000";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                
                      cntr <= "000100000001";
                elsif cntr ="000100000001" THEN
                      t1addb <= "10000001";
				      t2addb <= "10100001";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                
                
                      
				        zetain   <="00000100";
				      cntr <= "000100000010";
				elsif cntr ="000100000010" THEN
                      t1addb <= "10000010";
                      t2addb <= "10100010";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;      
                      
                      
                      
                
                      cntr <= "000100000011";
                elsif cntr ="000100000011" THEN
                      t1addb <= "10000011";
                      t2addb <= "10100011";
                      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100000100";
				elsif cntr ="000100000100" THEN
				      t1addb <= "10000100";
				      t2addb <= "10100100";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100000101";
				elsif cntr ="000100000101" THEN
				      t1addb <= "10000101";
				      t2addb <= "10100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100000110";
				elsif cntr ="000100000110" THEN
				      t1addb <= "10000110";      
				      t2addb <= "10100110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100000111";
				elsif cntr ="000100000111" THEN
				      t1addb <= "10000111";
				      t2addb <= "10100111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100001000";
				elsif cntr ="000100001000" THEN
				      t1addb <= "10001000";
				      t2addb <= "10101000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000100001001";
				elsif cntr ="000100001001" THEN
				      t1addb <= "10001001";
				      t2addb <= "10101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      cntr <= "000100001010";
				elsif cntr ="000100001010" THEN
				      t1addb <= "10001010";
				      t2addb <= "10101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100001011";
				elsif cntr ="000100001011" THEN
				      t1addb <= "10001011";
				      t2addb <= "10101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000100001100";
				elsif cntr ="000100001100" THEN
				      t1addb <= "10001100";
				      t2addb <= "10101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100001101";
				elsif cntr ="000100001101" THEN
				      t1addb <= "10001101";
				      t2addb <= "10101101";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100001110";
				elsif cntr ="000100001110" THEN
				      t1addb <= "10001110";
				      t2addb <= "10101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100001111";
				elsif cntr ="000100001111" THEN
				      t1addb <= "10001111";
                      t2addb <= "10101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010000";
				elsif cntr ="000100010000" THEN
				      t1addb <= "10010000";
				      t2addb <= "10110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010001";
                elsif cntr ="000100010001" THEN
				      t1addb <= "10010001";
				      t2addb <= "10110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010010";
				elsif cntr ="000100010010" THEN
				      t1addb <= "10010010";
				      t2addb <= "10110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000100010011";
				elsif cntr ="000100010011" THEN
				      t1addb <= "10010011";
				      t2addb <= "10110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010100";
				elsif cntr ="000100010100" THEN
				      t1addb <= "10010100";
				      t2addb <= "10110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010101";
				elsif cntr ="000100010101" THEN
				      t1addb <= "10010101";
				      t2addb <= "10110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010110";
				elsif cntr ="000100010110" THEN
				      t1addb <= "10010110";
				      t2addb <= "10110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100010111";
				elsif cntr ="000100010111" THEN
				      t1addb <= "10010111";
				      t2addb <= "10110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011000";
				elsif cntr ="000100011000" THEN
				      t1addb <= "10011000";
				      t2addb <= "10111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011001";
				elsif cntr ="000100011001" THEN
				      t1addb <= "10011001";
				      t2addb <= "10111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011010";
				elsif cntr ="000100011010" THEN
				      t1addb <= "10011010";
				      t2addb <= "10111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011011";
				elsif cntr ="000100011011" THEN
				      t1addb <= "10011011";
				      t2addb <= "10111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011100";
				elsif cntr ="000100011100" THEN
				      t1addb <= "10011100";
				      t2addb <= "10111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000100011101";
				elsif cntr ="000100011101" THEN
				      t1addb <= "10011101";
				      t2addb <= "10111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011110";
				elsif cntr ="000100011110" THEN
				      t1addb <= "10011110";
				      t2addb <= "10111110";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100011111";
				elsif cntr ="000100011111" THEN
				      t1addb <= "10011111";
				      t2addb <= "10111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100100000";
				elsif cntr ="000100100000" THEN
				      t1addb <= "10100000";
                      t2addb <= "10000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000100100001";
				elsif cntr ="000100100001" THEN
				      t1addb <= "10100001";
				      t2addb <= "10000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00000101";
				      cntr <= "000100100010";
                elsif cntr ="000100100010" THEN
				      t1addb <= "10100010";
				      t2addb <= "10000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100100011";
				elsif cntr ="000100100011" THEN
				      t1addb <= "10100011";
				      t2addb <= "10000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "000100100100";
				elsif cntr ="000100100100" THEN
				      t1addb <= "10100100";
				      t2addb <= "10000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100100101";
				elsif cntr ="000100100101" THEN
				      t1addb <= "10100101";
				      t2addb <= "10000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100100110";
				elsif cntr ="000100100110" THEN
				      t1addb <= "10100110";
				      t2addb <= "10000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100100111";
				elsif cntr ="000100100111" THEN
				      t1addb <= "10100111";
				      t2addb <= "10000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101000";
				elsif cntr ="000100101000" THEN
				      t1addb <= "10101000";
				      t2addb <= "10001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101001";
				elsif cntr ="000100101001" THEN
				      t1addb <= "10101001";
				      t2addb <= "10001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101010";
				elsif cntr ="000100101010" THEN
				      t1addb <= "10101010";
				      t2addb <= "10001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101011";
				elsif cntr ="000100101011" THEN
				      t1addb <= "10101011";
				      t2addb <= "10001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101100";
				elsif cntr ="000100101100" THEN
				      t1addb <= "10101100";
				      t2addb <= "10001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101101";
				elsif cntr ="000100101101" THEN
				      t1addb <= "10101101";
				      t2addb <= "10001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "000100101110";
				elsif cntr ="000100101110" THEN
				      t1addb <= "10101110";
				      t2addb <= "10001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100101111";
				elsif cntr ="000100101111" THEN
				      t1addb <= "10101111";
				      t2addb <= "10001111";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110000";
				elsif cntr ="000100110000" THEN
				      t1addb <= "10110000";
				      t2addb <= "10010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110001";
				elsif cntr ="000100110001" THEN
				      t1addb <= "10110001";
                      t2addb <= "10010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110010";
				elsif cntr ="000100110010" THEN
				      t1addb <= "10110010";
				      t2addb <= "10010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110011";
                elsif cntr ="000100110011" THEN
				      t1addb <= "10110011";
				      t2addb <= "10010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110100";
				elsif cntr ="000100110100" THEN
				      t1addb <= "10110100";
				      t2addb <= "10010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "000100110101";
				elsif cntr ="000100110101" THEN
				      t1addb <= "10110101";
				      t2addb <= "10010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110110";
				elsif cntr ="000100110110" THEN
				      t1addb <= "10110110";
				      t2addb <= "10010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100110111";
				elsif cntr ="000100110111" THEN
				      t1addb <= "10110111";
				      t2addb <= "10010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111000";
				elsif cntr ="000100111000" THEN
				      t1addb <= "10111000";
				      t2addb <= "10011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111001";
				elsif cntr ="000100111001" THEN
				      t1addb <= "10111001";
				      t2addb <= "10011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111010";
				elsif cntr ="000100111010" THEN
				      t1addb <= "10111010";
				      t2addb <= "10011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111011";
				elsif cntr ="000100111011" THEN
				      t1addb <= "10111011";
				      t2addb <= "10011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111100";
				elsif cntr ="000100111100" THEN
				      t1addb <= "10111100";
				      t2addb <= "10011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111101";
				elsif cntr ="000100111101" THEN
				      t1addb <= "10111101";
				      t2addb <= "10011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000100111110";
				elsif cntr ="000100111110" THEN
				      t1addb <= "10111110";
				      t2addb <= "10011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "000100111111";
				elsif cntr ="000100111111" THEN
				      t1addb <= "10111111";
				      t2addb <= "10011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101000000";
				elsif cntr ="000101000000" THEN
				      t1addb <= "11000000";
				      t2addb <= "11100000";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101000001";
				elsif cntr ="000101000001" THEN
				      t1addb <= "11000001";
				      t2addb <= "11100001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00000110";
				      cntr <= "000101000010";
				elsif cntr ="000101000010" THEN
				      t1addb <= "11000010";
                      t2addb <= "11100010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101000011";
				elsif cntr ="000101000011" THEN
				      t1addb <= "11000011";
				      t2addb <= "11100011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101000100";
                elsif cntr ="000101000100" THEN
				      t1addb <= "11000100";
				      t2addb <= "11100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101000101";
				elsif cntr ="000101000101" THEN
				      t1addb <= "11000101";
				      t2addb <= "11100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000101000110";
				elsif cntr ="000101000110" THEN
				      t1addb <= "11000110";
				      t2addb <= "11100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101000111";
				elsif cntr ="000101000111" THEN
				      t1addb <= "11000111";
				      t2addb <= "11100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001000";
				elsif cntr ="000101001000" THEN
				      t1addb <= "11001000";
				      t2addb <= "11101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001001";
				elsif cntr ="000101001001" THEN
				      t1addb <= "11001001";
				      t2addb <= "11101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001010";
				elsif cntr ="000101001010" THEN
				      t1addb <= "11001010";
				      t2addb <= "11101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001011";
				elsif cntr ="000101001011" THEN
				      t1addb <= "11001011";
				      t2addb <= "11101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001100";
				elsif cntr ="000101001100" THEN
				      t1addb <= "11001100";
				      t2addb <= "11101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001101";
				elsif cntr ="000101001101" THEN
				      t1addb <= "11001101";
				      t2addb <= "11101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001110";
				elsif cntr ="000101001110" THEN
				      t1addb <= "11001110";
				      t2addb <= "11101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101001111";
				elsif cntr ="000101001111" THEN
				      t1addb <= "11001111";
				      t2addb <= "11101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000101010000";
				elsif cntr ="000101010000" THEN
				      t1addb <= "11010000";
				      t2addb <= "11110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010001";
				elsif cntr ="000101010001" THEN
				      t1addb <= "11010001";
				      t2addb <= "11110001";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010010";
				elsif cntr ="000101010010" THEN
				      t1addb <= "11010010";
				      t2addb <= "11110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010011";
				elsif cntr ="000101010011" THEN
				      t1addb <= "11010011";
                      t2addb <= "11110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010100";
				elsif cntr ="000101010100" THEN
				      t1addb <= "11010100";
				      t2addb <= "11110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010101";
                elsif cntr ="000101010101" THEN
				      t1addb <= "11010101";
				      t2addb <= "11110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101010110";
				elsif cntr ="000101010110" THEN
				      t1addb <= "11010110";
				      t2addb <= "11110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000101010111";
				elsif cntr ="000101010111" THEN
				      t1addb <= "11010111";
				      t2addb <= "11110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011000";
				elsif cntr ="000101011000" THEN
				      t1addb <= "11011000";
				      t2addb <= "11111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011001";
				elsif cntr ="000101011001" THEN
				      t1addb <= "11011001";
				      t2addb <= "11111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011010";
				elsif cntr ="000101011010" THEN
				      t1addb <= "11011010";
				      t2addb <= "11111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011011";
				elsif cntr ="000101011011" THEN
				      t1addb <= "11011011";
				      t2addb <= "11111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011100";
				elsif cntr ="000101011100" THEN
				      t1addb <= "11011100";
				      t2addb <= "11111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011101";
				elsif cntr ="000101011101" THEN
				      t1addb <= "11011101";
				      t2addb <= "11111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011110";
				elsif cntr ="000101011110" THEN
				      t1addb <= "11011110";
				      t2addb <= "11111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101011111";
				elsif cntr ="000101011111" THEN
				      t1addb <= "11011111";
				      t2addb <= "11111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000101100000";
				elsif cntr ="000101100000" THEN
				      t1addb <= "11100000";
				      t2addb <= "11000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000101100001";
				elsif cntr ="000101100001" THEN
				      t1addb <= "11100001";
				      t2addb <= "11000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00000111";
				      cntr <= "000101100010";
				elsif cntr ="000101100010" THEN
				      t1addb <= "11100010";
				      t2addb <= "11000010";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101100011";
				elsif cntr ="000101100011" THEN
				      t1addb <= "11100011";
				      t2addb <= "11000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101100100";
				elsif cntr ="000101100100" THEN
				      t1addb <= "11100100";
                      t2addb <= "11000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101100101";
				elsif cntr ="000101100101" THEN
				      t1addb <= "11100101";
				      t2addb <= "11000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101100110";
                elsif cntr ="000101100110" THEN
				      t1addb <= "11100110";
				      t2addb <= "11000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101100111";
				elsif cntr ="000101100111" THEN
				      t1addb <= "11100111";
				      t2addb <= "11000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "000101101000";
				elsif cntr ="000101101000" THEN
				      t1addb <= "11101000";
				      t2addb <= "11001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101001";
				elsif cntr ="000101101001" THEN
				      t1addb <= "11101001";
				      t2addb <= "11001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101010";
				elsif cntr ="000101101010" THEN
				      t1addb <= "11101010";
				      t2addb <= "11001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101011";
				elsif cntr ="000101101011" THEN
				      t1addb <= "11101011";
				      t2addb <= "11001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101100";
				elsif cntr ="000101101100" THEN
				      t1addb <= "11101100";
				      t2addb <= "11001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101101";
				elsif cntr ="000101101101" THEN
				      t1addb <= "11101101";
				      t2addb <= "11001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101110";
				elsif cntr ="000101101110" THEN
				      t1addb <= "11101110";
				      t2addb <= "11001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101101111";
				elsif cntr ="000101101111" THEN
				      t1addb <= "11101111";
				      t2addb <= "11001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110000";
				elsif cntr ="000101110000" THEN
				      t1addb <= "11110000";
				      t2addb <= "11010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110001";
				elsif cntr ="000101110001" THEN
				      t1addb <= "11110001";
				      t2addb <= "11010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "000101110010";
				elsif cntr ="000101110010" THEN
				      t1addb <= "11110010";
				      t2addb <= "11010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110011";
				elsif cntr ="000101110011" THEN
				      t1addb <= "11110011";
				      t2addb <= "11010011";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110100";
				elsif cntr ="000101110100" THEN
				      t1addb <= "11110100";
				      t2addb <= "11010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110101";
				elsif cntr ="000101110101" THEN
				      t1addb <= "11110101";
                      t2addb <= "11010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110110";
				elsif cntr ="000101110110" THEN
				      t1addb <= "11110110";
				      t2addb <= "11010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101110111";
                elsif cntr ="000101110111" THEN
				      t1addb <= "11110111";
				      t2addb <= "11010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111000";
				elsif cntr ="000101111000" THEN
				      t1addb <= "11111000";
				      t2addb <= "11011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "000101111001";
				elsif cntr ="000101111001" THEN
				      t1addb <= "11111001";
				      t2addb <= "11011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111010";
				elsif cntr ="000101111010" THEN
				      t1addb <= "11111010";
				      t2addb <= "11011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111011";
				elsif cntr ="000101111011" THEN
				      t1addb <= "11111011";
				      t2addb <= "11011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111100";
				elsif cntr ="000101111100" THEN
				      t1addb <= "11111100";
				      t2addb <= "11011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111101";
				elsif cntr ="000101111101" THEN
				      t1addb <= "11111101";
				      t2addb <= "11011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111110";
				elsif cntr ="000101111110" THEN
				      t1addb <= "11111110";
				      t2addb <= "11011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000101111111";
				elsif cntr ="000101111111" THEN
				      t1addb <= "11111111";
				      t2addb <= "11011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110000000";
				elsif cntr ="000110000000" THEN
                      t1addb <= "00000000";
                      t2addb <= "00010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				      
				      
				      
				      cntr <= "000110000001";
				elsif cntr ="000110000001" THEN
                      t1addb <= "00000001";
                      t2addb <= "00010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				
				      
				        zetain   <="00001000";      
				      cntr <= "000110000010";
				elsif cntr ="000110000010" THEN
				      t1addb <= "00000010";
				      t2addb <= "00010010";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
                      
				            
				      cntr <= "000110000011";
				elsif cntr ="000110000011" THEN    
				      t1addb <= "00000011";
				      t2addb <= "00010011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
                
                      cntr <= "000110000100";
                elsif cntr ="000110000100" THEN
                      t1addb <= "00000100";
                      t2addb <= "00010100";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
                      
				      
				      
				
				      cntr <= "000110000101";     
				elsif cntr ="000110000101" THEN     
				      t1addb <= "00000101";
				      t2addb <= "00010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000110000110";         
				elsif cntr ="000110000110" THEN         
				      t1addb <= "00000110";
				      t2addb <= "00010110";
                      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000110000111";
				elsif cntr ="000110000111" THEN
				      t1addb <= "00000111";
				      t2addb <= "00010111";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				  
				      cntr <= "000110001000";  
				elsif cntr ="000110001000" THEN  
                      t1addb <= "00001000";
				      t2addb <= "00011000";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "000110001001";
				elsif cntr ="000110001001" THEN
				      t1addb <= "00001001";
				      t2addb <= "00011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
					  
				
				
				      
                      cntr <= "000110001010";
				elsif cntr ="000110001010" THEN
				      t1addb <= "00001010";
				      t2addb <= "00011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110001011";
				elsif cntr ="000110001011" THEN
				      t1addb <= "00001011";
				      t2addb <= "00011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110001100";
				elsif cntr ="000110001100" THEN
				      t1addb <= "00001100";
				      t2addb <= "00011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110001101";
				elsif cntr ="000110001101" THEN
				      t1addb <= "00001101";
				      t2addb <= "00011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110001110";
				elsif cntr ="000110001110" THEN
				      t1addb <= "00001110";
				      t2addb <= "00011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110001111";
				elsif cntr ="000110001111" THEN
				      t1addb <= "00001111";
                      t2addb <= "00011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110010000";
				elsif cntr ="000110010000" THEN
				      t1addb <= "00010000";
				      t2addb <= "00000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110010001";
				elsif cntr ="000110010001" THEN
				      t1addb <= "00010001";
				      t2addb <= "00000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00001001";
				      cntr <= "000110010010";
				elsif cntr ="000110010010" THEN
				      t1addb <= "00010010";
				      t2addb <= "00000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "000110010011";
				elsif cntr ="000110010011" THEN
				      t1addb <= "00010011";
				      t2addb <= "00000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
                      cntr <= "000110010100";
				elsif cntr ="000110010100" THEN
				      t1addb <= "00010100";
				      t2addb <= "00000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110010101";
				elsif cntr ="000110010101" THEN
				      t1addb <= "00010101";
				      t2addb <= "00000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110010110";
				elsif cntr ="000110010110" THEN
				      t1addb <= "00010110";
				      t2addb <= "00000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110010111";
				elsif cntr ="000110010111" THEN
				      t1addb <= "00010111";
				      t2addb <= "00000111";
                      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011000";
				elsif cntr ="000110011000" THEN
				      t1addb <= "00011000";
				      t2addb <= "00001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011001";
				elsif cntr ="000110011001" THEN
				      t1addb <= "00011001";
				      t2addb <= "00001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011010";
				elsif cntr ="000110011010" THEN
				      t1addb <= "00011010";
				      t2addb <= "00001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
                      
				      
				      cntr <= "000110011011";
				elsif cntr ="000110011011" THEN
				      t1addb <= "00011011";
				      t2addb <= "00001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011100";
                elsif cntr ="000110011100" THEN
				      t1addb <= "00011100";
				      t2addb <= "00001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011101";
				elsif cntr ="000110011101" THEN
				      t1addb <= "00011101";
				      t2addb <= "00001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011110";
				elsif cntr ="000110011110" THEN
				      t1addb <= "00011110";
				      t2addb <= "00001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110011111";
				elsif cntr ="000110011111" THEN
				      t1addb <= "00011111";
				      t2addb <= "00001111";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110100000";
				elsif cntr ="000110100000" THEN
				      t1addb <= "00100000";
				      t2addb <= "00110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110100001";
				elsif cntr ="000110100001" THEN
				      t1addb <= "00100001";
				      t2addb <= "00110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00001010";
				      cntr <= "000110100010";
				elsif cntr ="000110100010" THEN
				      t1addb <= "00100010";
				      t2addb <= "00110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110100011";
				elsif cntr ="000110100011" THEN
				      t1addb <= "00100011";
				      t2addb <= "00110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110100100";
				elsif cntr ="000110100100" THEN
                      t1addb <= "00100100";
				      t2addb <= "00110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110100101";
				elsif cntr ="000110100101" THEN
				      t1addb <= "00100101";
				      t2addb <= "00110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110100110";
				elsif cntr ="000110100110" THEN
				      t1addb <= "00100110";
				      t2addb <= "00110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110100111";
				elsif cntr ="000110100111" THEN
				      t1addb <= "00100111";
				      t2addb <= "00110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
                      
				      
				      
				      
				      cntr <= "000110101000";
				elsif cntr ="000110101000" THEN
				      t1addb <= "00101000";
				      t2addb <= "00111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000110101001";
				elsif cntr ="000110101001" THEN
				      t1addb <= "00101001";
				      t2addb <= "00111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101010";
				elsif cntr ="000110101010" THEN
				      t1addb <= "00101010";
				      t2addb <= "00111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101011";
				elsif cntr ="000110101011" THEN
				      t1addb <= "00101011";
				      t2addb <= "00111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101100";
				elsif cntr ="000110101100" THEN
				      t1addb <= "00101100";
                      t2addb <= "00111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101101";
				elsif cntr ="000110101101" THEN
				      t1addb <= "00101101";
				      t2addb <= "00111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101110";
				elsif cntr ="000110101110" THEN
				      t1addb <= "00101110";
				      t2addb <= "00111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000110101111";
				elsif cntr ="000110101111" THEN
				      t1addb <= "00101111";
				      t2addb <= "00111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000110110000";
				elsif cntr ="000110110000" THEN
				      t1addb <= "00110000";
				      t2addb <= "00100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
                      cntr <= "000110110001";
				elsif cntr ="000110110001" THEN
				      t1addb <= "00110001";
				      t2addb <= "00100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00001011";
				      cntr <= "000110110010";
				elsif cntr ="000110110010" THEN
				      t1addb <= "00110010";
				      t2addb <= "00100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110110011";
				elsif cntr ="000110110011" THEN
				      t1addb <= "00110011";
				      t2addb <= "00100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110110100";
				elsif cntr ="000110110100" THEN
				      t1addb <= "00110100";
				      t2addb <= "00100100";
                      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110110101";
				elsif cntr ="000110110101" THEN
				      t1addb <= "00110101";
				      t2addb <= "00100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110110110";
				elsif cntr ="000110110110" THEN
				      t1addb <= "00110110";
				      t2addb <= "00100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110110111";
				elsif cntr ="000110110111" THEN
				      t1addb <= "00110111";
				      t2addb <= "00100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
                      
				      
				      cntr <= "000110111000";
				elsif cntr ="000110111000" THEN
				      t1addb <= "00111000";
				      t2addb <= "00101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111001";
                elsif cntr ="000110111001" THEN
				      t1addb <= "00111001";
				      t2addb <= "00101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111010";
				elsif cntr ="000110111010" THEN
				      t1addb <= "00111010";
				      t2addb <= "00101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111011";
				elsif cntr ="000110111011" THEN
				      t1addb <= "00111011";
				      t2addb <= "00101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111100";
				elsif cntr ="000110111100" THEN
				      t1addb <= "00111100";
				      t2addb <= "00101100";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111101";
				elsif cntr ="000110111101" THEN
				      t1addb <= "00111101";
				      t2addb <= "00101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111110";
				elsif cntr ="000110111110" THEN
				      t1addb <= "00111110";
				      t2addb <= "00101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000110111111";
				elsif cntr ="000110111111" THEN
				      t1addb <= "00111111";
				      t2addb <= "00101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111000000";
				elsif cntr ="000111000000" THEN
				      t1addb <= "01000000";
				      t2addb <= "01010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111000001";
				elsif cntr ="000111000001" THEN
                      t1addb <= "01000001";
				      t2addb <= "01010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00001100";
				      cntr <= "000111000010";
				elsif cntr ="000111000010" THEN
				      t1addb <= "01000010";
				      t2addb <= "01010010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111000011";
				elsif cntr ="000111000011" THEN
				      t1addb <= "01000011";
				      t2addb <= "01010011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111000100";
				elsif cntr ="000111000100" THEN
				      t1addb <= "01000100";
				      t2addb <= "01010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
                      
				      
				      
				      
				      cntr <= "000111000101";
				elsif cntr ="000111000101" THEN
				      t1addb <= "01000101";
				      t2addb <= "01010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000111000110";
				elsif cntr ="000111000110" THEN
				      t1addb <= "01000110";
				      t2addb <= "01010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111000111";
				elsif cntr ="000111000111" THEN
				      t1addb <= "01000111";
				      t2addb <= "01010111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001000";
				elsif cntr ="000111001000" THEN
				      t1addb <= "01001000";
				      t2addb <= "01011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001001";
				elsif cntr ="000111001001" THEN
				      t1addb <= "01001001";
                      t2addb <= "01011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001010";
				elsif cntr ="000111001010" THEN
				      t1addb <= "01001010";
				      t2addb <= "01011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001011";
				elsif cntr ="000111001011" THEN
				      t1addb <= "01001011";
				      t2addb <= "01011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001100";
				elsif cntr ="000111001100" THEN
				      t1addb <= "01001100";
				      t2addb <= "01011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000111001101";
				elsif cntr ="000111001101" THEN
				      t1addb <= "01001101";
				      t2addb <= "01011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
                      cntr <= "000111001110";
				elsif cntr ="000111001110" THEN
				      t1addb <= "01001110";
				      t2addb <= "01011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111001111";
				elsif cntr ="000111001111" THEN
				      t1addb <= "01001111";
				      t2addb <= "01011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111010000";
				elsif cntr ="000111010000" THEN
				      t1addb <= "01010000";
				      t2addb <= "01000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111010001";
				elsif cntr ="000111010001" THEN
				      t1addb <= "01010001";
				      t2addb <= "01000001";
                      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00001101";
				      cntr <= "000111010010";
				elsif cntr ="000111010010" THEN
				      t1addb <= "01010010";
				      t2addb <= "01000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111010011";
				elsif cntr ="000111010011" THEN
				      t1addb <= "01010011";
				      t2addb <= "01000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111010100";
				elsif cntr ="000111010100" THEN
				      t1addb <= "01010100";
				      t2addb <= "01000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
                      
				      
				      cntr <= "000111010101";
				elsif cntr ="000111010101" THEN
				      t1addb <= "01010101";
				      t2addb <= "01000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111010110";
                elsif cntr ="000111010110" THEN
				      t1addb <= "01010110";
				      t2addb <= "01000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111010111";
				elsif cntr ="000111010111" THEN
				      t1addb <= "01010111";
				      t2addb <= "01000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011000";
				elsif cntr ="000111011000" THEN
				      t1addb <= "01011000";
				      t2addb <= "01001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011001";
				elsif cntr ="000111011001" THEN
				      t1addb <= "01011001";
				      t2addb <= "01001001";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011010";
				elsif cntr ="000111011010" THEN
				      t1addb <= "01011010";
				      t2addb <= "01001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011011";
				elsif cntr ="000111011011" THEN
				      t1addb <= "01011011";
				      t2addb <= "01001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011100";
				elsif cntr ="000111011100" THEN
				      t1addb <= "01011100";
				      t2addb <= "01001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011101";
				elsif cntr ="000111011101" THEN
				      t1addb <= "01011101";
				      t2addb <= "01001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011110";
				elsif cntr ="000111011110" THEN
                      t1addb <= "01011110";
				      t2addb <= "01001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111011111";
				elsif cntr ="000111011111" THEN
				      t1addb <= "01011111";
				      t2addb <= "01001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111100000";
				elsif cntr ="000111100000" THEN
				      t1addb <= "01100000";
				      t2addb <= "01110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111100001";
				elsif cntr ="000111100001" THEN
				      t1addb <= "01100001";
				      t2addb <= "01110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
                      
				      
				      
				        zetain   <="00001110";
				      cntr <= "000111100010";
				elsif cntr ="000111100010" THEN
				      t1addb <= "01100010";
				      t2addb <= "01110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
                      
				      cntr <= "000111100011";
				elsif cntr ="000111100011" THEN
				      t1addb <= "01100011";
				      t2addb <= "01110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111100100";
				elsif cntr ="000111100100" THEN
				      t1addb <= "01100100";
				      t2addb <= "01110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111100101";
				elsif cntr ="000111100101" THEN
				      t1addb <= "01100101";
				      t2addb <= "01110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111100110";
				elsif cntr ="000111100110" THEN
				      t1addb <= "01100110";
                      t2addb <= "01110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111100111";
				elsif cntr ="000111100111" THEN
				      t1addb <= "01100111";
				      t2addb <= "01110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101000";
				elsif cntr ="000111101000" THEN
				      t1addb <= "01101000";
				      t2addb <= "01111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101001";
				elsif cntr ="000111101001" THEN
				      t1addb <= "01101001";
				      t2addb <= "01111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "000111101010";
				elsif cntr ="000111101010" THEN
				      t1addb <= "01101010";
				      t2addb <= "01111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
                      cntr <= "000111101011";
				elsif cntr ="000111101011" THEN
				      t1addb <= "01101011";
				      t2addb <= "01111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101100";
				elsif cntr ="000111101100" THEN
				      t1addb <= "01101100";
				      t2addb <= "01111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101101";
				elsif cntr ="000111101101" THEN
				      t1addb <= "01101101";
				      t2addb <= "01111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101110";
				elsif cntr ="000111101110" THEN
				      t1addb <= "01101110";
				      t2addb <= "01111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111101111";
				elsif cntr ="000111101111" THEN
				      t1addb <= "01101111";
				      t2addb <= "01111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111110000";
				elsif cntr ="000111110000" THEN
				      t1addb <= "01110000";
				      t2addb <= "01100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "000111110001";
				elsif cntr ="000111110001" THEN
				      t1addb <= "01110001";
				      t2addb <= "01100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00001111";
				      cntr <= "000111110010";
				elsif cntr ="000111110010" THEN
				      t1addb <= "01110010";
				      t2addb <= "01100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111110011";
				elsif cntr ="000111110011" THEN
				      t1addb <= "01110011";
				      t2addb <= "01100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111110100";
				elsif cntr ="000111110100" THEN
				      t1addb <= "01110100";
				      t2addb <= "01100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "000111110101";
				elsif cntr ="000111110101" THEN
				      t1addb <= "01110101";
				      t2addb <= "01100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111110110";
				elsif cntr ="000111110110" THEN
				      t1addb <= "01110110";
				      t2addb <= "01100110";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111110111";
				elsif cntr ="000111110111" THEN
				      t1addb <= "01110111";
				      t2addb <= "01100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111000";
				elsif cntr ="000111111000" THEN
				      t1addb <= "01111000";
				      t2addb <= "01101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111001";
				elsif cntr ="000111111001" THEN
				      t1addb <= "01111001";
				      t2addb <= "01101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111010";
				elsif cntr ="000111111010" THEN
				      t1addb <= "01111010";
				      t2addb <= "01101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111011";
				elsif cntr ="000111111011" THEN
				      t1addb <= "01111011";
				      t2addb <= "01101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111100";
				elsif cntr ="000111111100" THEN
				      t1addb <= "01111100";
				      t2addb <= "01101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
                      
				      
				      cntr <= "000111111101";
				elsif cntr ="000111111101" THEN
				      t1addb <= "01111101";
				      t2addb <= "01101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111110";
				elsif cntr ="000111111110" THEN
				      t1addb <= "01111110";
				      t2addb <= "01101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "000111111111";
				elsif cntr ="000111111111" THEN
				      t1addb <= "01111111";
				      t2addb <= "01101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000000000";
				elsif cntr ="001000000000" THEN
				      t1addb <= "10000000";
				      t2addb <= "10001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000000001";
				elsif cntr ="001000000001" THEN
				      t1addb <= "10000001";
				      t2addb <= "10001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				      
				      
				        zetain   <="00010000";      
				      cntr <= "001000000010";
				elsif cntr ="001000000010" THEN
				      t1addb <= "10000010";
				      t2addb <= "10001010";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				      cntr <= "001000000011";
				elsif cntr ="001000000011" THEN
				      t1addb <= "10000011";
				      t2addb <= "10001011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				                  
				      cntr <= "001000000100";
				elsif cntr ="001000000100" THEN
				      t1addb <= "10000100";
				      t2addb <= "10001100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				      cntr <= "001000000101";
				elsif cntr ="001000000101" THEN
				      t1addb <= "10000101";
				      t2addb <= "10001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;      
				      
				      
				      
                                              
				      cntr <= "001000000110";
				elsif cntr ="001000000110" THEN
				      t1addb <= "10000110";
				      t2addb <= "10001110";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "001000000111";
				elsif cntr ="001000000111" THEN
				      t1addb <= "10000111";      
				      t2addb <= "10001111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				    
				      cntr <= "001000001000";     
				elsif cntr ="001000001000" THEN     
				      t1addb <= "10001000";
				      t2addb <= "10000000";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "001000001001";
				elsif cntr ="001000001001" THEN
				      t1addb <= "10001001";
				      t2addb <= "10000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
					  
				
				
				        zetain   <="00010001";
				      cntr <= "001000001010";
				elsif cntr ="001000001010" THEN
				      t1addb <= "10001010";
				      t2addb <= "10000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000001011";
				elsif cntr ="001000001011" THEN
				      t1addb <= "10001011";
				      t2addb <= "10000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000001100";
				elsif cntr ="001000001100" THEN
                      t1addb <= "10001100";
				      t2addb <= "10000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000001101";
				elsif cntr ="001000001101" THEN
				      t1addb <= "10001101";
				      t2addb <= "10000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
                      cntr <= "001000001110";
				elsif cntr ="001000001110" THEN
				      t1addb <= "10001110";
				      t2addb <= "10000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000001111";
				elsif cntr ="001000001111" THEN
				      t1addb <= "10001111";
				      t2addb <= "10000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000010000";
				elsif cntr ="001000010000" THEN
				      t1addb <= "10010000";
				      t2addb <= "10011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000010001";
				elsif cntr ="001000010001" THEN
				      t1addb <= "10010001";
				      t2addb <= "10011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00010010";
				      cntr <= "001000010010";
				elsif cntr ="001000010010" THEN
				      t1addb <= "10010010";
				      t2addb <= "10011010";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000010011";
				elsif cntr ="001000010011" THEN
				      t1addb <= "10010011";
				      t2addb <= "10011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000010100";
				elsif cntr ="001000010100" THEN
				      t1addb <= "10010100";
                      t2addb <= "10011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000010101";
				elsif cntr ="001000010101" THEN
				      t1addb <= "10010101";
				      t2addb <= "10011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000010110";
                elsif cntr ="001000010110" THEN
				      t1addb <= "10010110";
				      t2addb <= "10011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000010111";
				elsif cntr ="001000010111" THEN
				      t1addb <= "10010111";
				      t2addb <= "10011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000011000";
				elsif cntr ="001000011000" THEN
				      t1addb <= "10011000";
				      t2addb <= "10010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
                      
				      
				      cntr <= "001000011001";
				elsif cntr ="001000011001" THEN
				      t1addb <= "10011001";
				      t2addb <= "10010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00010011";
				      cntr <= "001000011010";
				elsif cntr ="001000011010" THEN
				      t1addb <= "10011010";
				      t2addb <= "10010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
                      
				      
				      
				      
				      cntr <= "001000011011";
				elsif cntr ="001000011011" THEN
				      t1addb <= "10011011";
				      t2addb <= "10010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000011100";
				elsif cntr ="001000011100" THEN
				      t1addb <= "10011100";
				      t2addb <= "10010100";
                      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000011101";
				elsif cntr ="001000011101" THEN
				      t1addb <= "10011101";
				      t2addb <= "10010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000011110";
				elsif cntr ="001000011110" THEN
				      t1addb <= "10011110";
				      t2addb <= "10010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000011111";
				elsif cntr ="001000011111" THEN
				      t1addb <= "10011111";
				      t2addb <= "10010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000100000";
				elsif cntr ="001000100000" THEN
				      t1addb <= "10100000";
				      t2addb <= "10101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000100001";
				elsif cntr ="001000100001" THEN
				      t1addb <= "10100001";
				      t2addb <= "10101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00010100";
				      cntr <= "001000100010";
				elsif cntr ="001000100010" THEN
				      t1addb <= "10100010";
				      t2addb <= "10101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "001000100011";
				elsif cntr ="001000100011" THEN
				      t1addb <= "10100011";
				      t2addb <= "10101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000100100";
				elsif cntr ="001000100100" THEN
				      t1addb <= "10100100";
				      t2addb <= "10101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000100101";
				elsif cntr ="001000100101" THEN
				      t1addb <= "10100101";
				      t2addb <= "10101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000100110";
				elsif cntr ="001000100110" THEN
				      t1addb <= "10100110";
				      t2addb <= "10101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000100111";
				elsif cntr ="001000100111" THEN
				      t1addb <= "10100111";
				      t2addb <= "10101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000101000";
				elsif cntr ="001000101000" THEN
				      t1addb <= "10101000";
				      t2addb <= "10100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000101001";
				elsif cntr ="001000101001" THEN
				      t1addb <= "10101001";
				      t2addb <= "10100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00010101";
				      cntr <= "001000101010";
				elsif cntr ="001000101010" THEN
				      t1addb <= "10101010";
				      t2addb <= "10100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "001000101011";
				elsif cntr ="001000101011" THEN
				      t1addb <= "10101011";
				      t2addb <= "10100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000101100";
				elsif cntr ="001000101100" THEN
				      t1addb <= "10101100";
				      t2addb <= "10100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000101101";
				elsif cntr ="001000101101" THEN
				      t1addb <= "10101101";
				      t2addb <= "10100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000101110";
				elsif cntr ="001000101110" THEN
				      t1addb <= "10101110";
				      t2addb <= "10100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000101111";
				elsif cntr ="001000101111" THEN
				      t1addb <= "10101111";
				      t2addb <= "10100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000110000";
				elsif cntr ="001000110000" THEN
				      t1addb <= "10110000";
				      t2addb <= "10111000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000110001";
				elsif cntr ="001000110001" THEN
                      t1addb <= "10110001";
				      t2addb <= "10111001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00010110";
				      cntr <= "001000110010";
				elsif cntr ="001000110010" THEN
				      t1addb <= "10110010";
				      t2addb <= "10111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
                      cntr <= "001000110011";
				elsif cntr ="001000110011" THEN
				      t1addb <= "10110011";
				      t2addb <= "10111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000110100";
				elsif cntr ="001000110100" THEN
				      t1addb <= "10110100";
				      t2addb <= "10111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000110101";
				elsif cntr ="001000110101" THEN
				      t1addb <= "10110101";
				      t2addb <= "10111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000110110";
				elsif cntr ="001000110110" THEN
				      t1addb <= "10110110";
				      t2addb <= "10111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000110111";
				elsif cntr ="001000110111" THEN
				      t1addb <= "10110111";
				      t2addb <= "10111111";
				      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000111000";
				elsif cntr ="001000111000" THEN
				      t1addb <= "10111000";
				      t2addb <= "10110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001000111001";
				elsif cntr ="001000111001" THEN
				      t1addb <= "10111001";
                      t2addb <= "10110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00010111";
				      cntr <= "001000111010";
				elsif cntr ="001000111010" THEN
				      t1addb <= "10111010";
				      t2addb <= "10110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000111011";
                elsif cntr ="001000111011" THEN
				      t1addb <= "10111011";
				      t2addb <= "10110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000111100";
				elsif cntr ="001000111100" THEN
				      t1addb <= "10111100";
				      t2addb <= "10110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000111101";
				elsif cntr ="001000111101" THEN
				      t1addb <= "10111101";
				      t2addb <= "10110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
                      
				      
				      cntr <= "001000111110";
				elsif cntr ="001000111110" THEN
				      t1addb <= "10111110";
				      t2addb <= "10110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001000111111";
				elsif cntr ="001000111111" THEN
				      t1addb <= "10111111";
				      t2addb <= "10110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
                      
				      
				      
				      
				      cntr <= "001001000000";
				elsif cntr ="001001000000" THEN
				      t1addb <= "11000000";
				      t2addb <= "11001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001000001";
				elsif cntr ="001001000001" THEN
				      t1addb <= "11000001";
				      t2addb <= "11001001";
                      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00011000";
				      cntr <= "001001000010";
				elsif cntr ="001001000010" THEN
				      t1addb <= "11000010";
				      t2addb <= "11001010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001000011";
				elsif cntr ="001001000011" THEN
				      t1addb <= "11000011";
				      t2addb <= "11001011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001000100";
				elsif cntr ="001001000100" THEN
				      t1addb <= "11000100";
				      t2addb <= "11001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001000101";
				elsif cntr ="001001000101" THEN
				      t1addb <= "11000101";
				      t2addb <= "11001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001000110";
				elsif cntr ="001001000110" THEN
				      t1addb <= "11000110";
				      t2addb <= "11001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001000111";
				elsif cntr ="001001000111" THEN
				      t1addb <= "11000111";
				      t2addb <= "11001111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
                      
				      
				      
				      cntr <= "001001001000";
				elsif cntr ="001001001000" THEN
				      t1addb <= "11001000";
				      t2addb <= "11000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001001001";
				elsif cntr ="001001001001" THEN
				      t1addb <= "11001001";
				      t2addb <= "11000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00011001";
				      cntr <= "001001001010";
				elsif cntr ="001001001010" THEN
				      t1addb <= "11001010";
				      t2addb <= "11000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001001011";
				elsif cntr ="001001001011" THEN
				      t1addb <= "11001011";
				      t2addb <= "11000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001001100";
				elsif cntr ="001001001100" THEN
				      t1addb <= "11001100";
				      t2addb <= "11000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001001101";
				elsif cntr ="001001001101" THEN
				      t1addb <= "11001101";
				      t2addb <= "11000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001001110";
				elsif cntr ="001001001110" THEN
				      t1addb <= "11001110";
				      t2addb <= "11000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001001111";
				elsif cntr ="001001001111" THEN
				      t1addb <= "11001111";
				      t2addb <= "11000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
                      
				      cntr <= "001001010000";
				elsif cntr ="001001010000" THEN
				      t1addb <= "11010000";
				      t2addb <= "11011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001010001";
				elsif cntr ="001001010001" THEN
				      t1addb <= "11010001";
				      t2addb <= "11011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00011010";
				      cntr <= "001001010010";
				elsif cntr ="001001010010" THEN
				      t1addb <= "11010010";
				      t2addb <= "11011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001010011";
				elsif cntr ="001001010011" THEN
				      t1addb <= "11010011";
				      t2addb <= "11011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001010100";
				elsif cntr ="001001010100" THEN
				      t1addb <= "11010100";
				      t2addb <= "11011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001010101";
				elsif cntr ="001001010101" THEN
				      t1addb <= "11010101";
				      t2addb <= "11011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001010110";
				elsif cntr ="001001010110" THEN
                      t1addb <= "11010110";
				      t2addb <= "11011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001010111";
				elsif cntr ="001001010111" THEN
				      t1addb <= "11010111";
				      t2addb <= "11011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
                      cntr <= "001001011000";
				elsif cntr ="001001011000" THEN
				      t1addb <= "11011000";
				      t2addb <= "11010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001011001";
				elsif cntr ="001001011001" THEN
				      t1addb <= "11011001";
				      t2addb <= "11010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00011011";
				      cntr <= "001001011010";
				elsif cntr ="001001011010" THEN
				      t1addb <= "11011010";
				      t2addb <= "11010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001011011";
				elsif cntr ="001001011011" THEN
				      t1addb <= "11011011";
				      t2addb <= "11010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001011100";
				elsif cntr ="001001011100" THEN
				      t1addb <= "11011100";
				      t2addb <= "11010100";
				      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001011101";
				elsif cntr ="001001011101" THEN
				      t1addb <= "11011101";
				      t2addb <= "11010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001011110";
				elsif cntr ="001001011110" THEN
				      t1addb <= "11011110";
                      t2addb <= "11010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001011111";
				elsif cntr ="001001011111" THEN
				      t1addb <= "11011111";
				      t2addb <= "11010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001100000";
                elsif cntr ="001001100000" THEN
				      t1addb <= "11100000";
				      t2addb <= "11101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001100001";
				elsif cntr ="001001100001" THEN
				      t1addb <= "11100001";
				      t2addb <= "11101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00011100";
				      cntr <= "001001100010";
				elsif cntr ="001001100010" THEN
				      t1addb <= "11100010";
				      t2addb <= "11101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
                      
				      
				      cntr <= "001001100011";
				elsif cntr ="001001100011" THEN
				      t1addb <= "11100011";
				      t2addb <= "11101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001100100";
				elsif cntr ="001001100100" THEN
				      t1addb <= "11100100";
				      t2addb <= "11101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
                      
				      
				      
				      
				      cntr <= "001001100101";
				elsif cntr ="001001100101" THEN
				      t1addb <= "11100101";
				      t2addb <= "11101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001100110";
				elsif cntr ="001001100110" THEN
				      t1addb <= "11100110";
				      t2addb <= "11101110";
                      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001100111";
				elsif cntr ="001001100111" THEN
				      t1addb <= "11100111";
				      t2addb <= "11101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001101000";
				elsif cntr ="001001101000" THEN
				      t1addb <= "11101000";
				      t2addb <= "11100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001101001";
				elsif cntr ="001001101001" THEN
				      t1addb <= "11101001";
				      t2addb <= "11100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00011101";
				      cntr <= "001001101010";
				elsif cntr ="001001101010" THEN
				      t1addb <= "11101010";
				      t2addb <= "11100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001101011";
				elsif cntr ="001001101011" THEN
				      t1addb <= "11101011";
				      t2addb <= "11100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001101100";
				elsif cntr ="001001101100" THEN
				      t1addb <= "11101100";
				      t2addb <= "11100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
                      
				      
				      
				      cntr <= "001001101101";
				elsif cntr ="001001101101" THEN
				      t1addb <= "11101101";
				      t2addb <= "11100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001101110";
				elsif cntr ="001001101110" THEN
				      t1addb <= "11101110";
				      t2addb <= "11100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001101111";
				elsif cntr ="001001101111" THEN
				      t1addb <= "11101111";
				      t2addb <= "11100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001110000";
				elsif cntr ="001001110000" THEN
				      t1addb <= "11110000";
				      t2addb <= "11111000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001110001";
				elsif cntr ="001001110001" THEN
				      t1addb <= "11110001";
				      t2addb <= "11111001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				        zetain   <="00011110";
				      cntr <= "001001110010";
				elsif cntr ="001001110010" THEN
				      t1addb <= "11110010";
				      t2addb <= "11111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001110011";
				elsif cntr ="001001110011" THEN
				      t1addb <= "11110011";
				      t2addb <= "11111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001110100";
				elsif cntr ="001001110100" THEN
				      t1addb <= "11110100";
				      t2addb <= "11111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
                      
				      
				      cntr <= "001001110101";
				elsif cntr ="001001110101" THEN
				      t1addb <= "11110101";
				      t2addb <= "11111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001110110";
				elsif cntr ="001001110110" THEN
				      t1addb <= "11110110";
				      t2addb <= "11111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
                      
				      
				      
				      
				      cntr <= "001001110111";
				elsif cntr ="001001110111" THEN
				      t1addb <= "11110111";
				      t2addb <= "11111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001111000";
				elsif cntr ="001001111000" THEN
				      t1addb <= "11111000";
				      t2addb <= "11110000";
                      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      cntr <= "001001111001";
				elsif cntr ="001001111001" THEN
				      t1addb <= "11111001";
				      t2addb <= "11110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				        zetain   <="00011111";
				      cntr <= "001001111010";
				elsif cntr ="001001111010" THEN
                      t1addb <= "11111010";
				      t2addb <= "11110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001111011";
				elsif cntr ="001001111011" THEN
				      t1addb <= "11111011";
				      t2addb <= "11110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
                      cntr <= "001001111100";
				elsif cntr ="001001111100" THEN
				      t1addb <= "11111100";
				      t2addb <= "11110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001111101";
				elsif cntr ="001001111101" THEN
				      t1addb <= "11111101";
				      t2addb <= "11110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001111110";
				elsif cntr ="001001111110" THEN
				      t1addb <= "11111110";
				      t2addb <= "11110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001001111111";
				elsif cntr ="001001111111" THEN
				      t1addb <= "11111111";
				      t2addb <= "11110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      cntr <= "001010000000";
				elsif cntr ="001010000000" THEN
				      t1addb <= "00000000";
				      t2addb <= "00000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				      
				      
				      
				      cntr <= "001010000001";
				elsif cntr ="001010000001" THEN
				      t1addb <= "00000001";
				      t2addb <= "00000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				      
				      
				        zetain   <="00100000";
				      cntr <= "001010000010";
				elsif cntr ="001010000010" THEN
				      t1addb <= "00000010";
				      t2addb <= "00000110";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				
				      cntr <= "001010000011";
				elsif cntr ="001010000011" THEN 
				      t1addb <= "00000011";
				      t2addb <= "00000111";
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
                                  
                      cntr <= "001010000100";
                elsif cntr ="001010000100" THEN
                      t1addb <= "00000100";
                      t2addb <= "00000000";
                      bfrjin     <= t1doutb;      
                      bfrjplin <= t2doutb;      
                      
                      
                      
                
                      cntr <= "001010000101";
                elsif cntr ="001010000101" THEN
                      t1addb <= "00000101";
                      t2addb <= "00000001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;      
                      
                      
                      
                        zetain   <="00100001";
                      cntr <= "001010000110";
                elsif cntr ="001010000110" THEN
                      t1addb <= "00000110";
                      t2addb <= "00000010";
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      
                      
                      
                
                      cntr <= "001010000111";
                elsif cntr ="001010000111" THEN
                      t1addb <= "00000111";
                      t2addb <= "00000011";
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      
                      
                      
                
                      cntr <= "001010001000";
                elsif cntr ="001010001000" THEN
                      t1addb <= "00001000";
                      t2addb <= "00001100";
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      
                      
                      
                
                      cntr <= "001010001001";
                elsif cntr ="001010001001" THEN
                      t1addb <= "00001001";
                      t2addb <= "00001101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      											
                
                
                        zetain   <="00100010";
                      cntr <= "001010001010";
                elsif cntr ="001010001010" THEN
                      t1addb <= "00001010";
                      t2addb <= "00001110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010001011";
                elsif cntr ="001010001011" THEN
                      t1addb <= "00001011";
                      t2addb <= "00001111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010001100";
                elsif cntr ="001010001100" THEN
                      t1addb <= "00001100";
                      t2addb <= "00001000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010001101";
                elsif cntr ="001010001101" THEN
                      t1addb <= "00001101";
                      t2addb <= "00001001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00100011";
                      cntr <= "001010001110";
                elsif cntr ="001010001110" THEN
                      t1addb <= "00001110";
                      t2addb <= "00001010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010001111";
                elsif cntr ="001010001111" THEN
                      t1addb <= "00001111";
                      t2addb <= "00001011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010010000";
                elsif cntr ="001010010000" THEN
                      t1addb <= "00010000";
                      t2addb <= "00010100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010010001";
                elsif cntr ="001010010001" THEN
                      t1addb <= "00010001";
                      t2addb <= "00010101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00100100";
                      cntr <= "001010010010";
                elsif cntr ="001010010010" THEN
                      t1addb <= "00010010";
                      t2addb <= "00010110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010010011";
                elsif cntr ="001010010011" THEN
                      t1addb <= "00010011";
                      t2addb <= "00010111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010010100";
                elsif cntr ="001010010100" THEN
                      t1addb <= "00010100";
                      t2addb <= "00010000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010010101";
                elsif cntr ="001010010101" THEN
                      t1addb <= "00010101";
                      t2addb <= "00010001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00100101";
                      cntr <= "001010010110";
                elsif cntr ="001010010110" THEN
                      t1addb <= "00010110";
                      t2addb <= "00010010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010010111";
                elsif cntr ="001010010111" THEN
                      t1addb <= "00010111";
                      t2addb <= "00010011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010011000";
                elsif cntr ="001010011000" THEN
                      t1addb <= "00011000";
                      t2addb <= "00011100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010011001";
                elsif cntr ="001010011001" THEN
                      t1addb <= "00011001";
                      t2addb <= "00011101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00100110";
                      cntr <= "001010011010";
                elsif cntr ="001010011010" THEN
                      t1addb <= "00011010";
                      t2addb <= "00011110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010011011";
                elsif cntr ="001010011011" THEN
                      t1addb <= "00011011";
                      t2addb <= "00011111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010011100";
                elsif cntr ="001010011100" THEN
                      t1addb <= "00011100";
                      t2addb <= "00011000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010011101";
                elsif cntr ="001010011101" THEN
                      t1addb <= "00011101";
                      t2addb <= "00011001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00100111";
                      cntr <= "001010011110";
                elsif cntr ="001010011110" THEN
                      t1addb <= "00011110";
                      t2addb <= "00011010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010011111";
                elsif cntr ="001010011111" THEN
                      t1addb <= "00011111";
                      t2addb <= "00011011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010100000";
                elsif cntr ="001010100000" THEN
                      t1addb <= "00100000";
                      t2addb <= "00100100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010100001";
                elsif cntr ="001010100001" THEN
                      t1addb <= "00100001";
                      t2addb <= "00100101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00101000";
                      cntr <= "001010100010";
                elsif cntr ="001010100010" THEN
                      t1addb <= "00100010";
                      t2addb <= "00100110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010100011";
                elsif cntr ="001010100011" THEN
                      t1addb <= "00100011";
                      t2addb <= "00100111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010100100";
                elsif cntr ="001010100100" THEN
                      t1addb <= "00100100";
                      t2addb <= "00100000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010100101";
                elsif cntr ="001010100101" THEN
                      t1addb <= "00100101";
                      t2addb <= "00100001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00101001";
                      cntr <= "001010100110";
                elsif cntr ="001010100110" THEN
                      t1addb <= "00100110";
                      t2addb <= "00100010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010100111";
                elsif cntr ="001010100111" THEN
                      t1addb <= "00100111";
                      t2addb <= "00100011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010101000";
                elsif cntr ="001010101000" THEN
                      t1addb <= "00101000";
                      t2addb <= "00101100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010101001";
                elsif cntr ="001010101001" THEN
                      t1addb <= "00101001";
                      t2addb <= "00101101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00101010";
                      cntr <= "001010101010";
                elsif cntr ="001010101010" THEN
                      t1addb <= "00101010";
                      t2addb <= "00101110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010101011";
                elsif cntr ="001010101011" THEN
                      t1addb <= "00101011";
                      t2addb <= "00101111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010101100";
                elsif cntr ="001010101100" THEN
                      t1addb <= "00101100";
                      t2addb <= "00101000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010101101";
                elsif cntr ="001010101101" THEN
                      t1addb <= "00101101";
                      t2addb <= "00101001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00101011";
                      cntr <= "001010101110";
                elsif cntr ="001010101110" THEN
                      t1addb <= "00101110";
                      t2addb <= "00101010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010101111";
                elsif cntr ="001010101111" THEN
                      t1addb <= "00101111";
                      t2addb <= "00101011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010110000";
                elsif cntr ="001010110000" THEN
                      t1addb <= "00110000";
                      t2addb <= "00110100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010110001";
                elsif cntr ="001010110001" THEN
                      t1addb <= "00110001";
                      t2addb <= "00110101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00101100";
                      cntr <= "001010110010";
                elsif cntr ="001010110010" THEN
                      t1addb <= "00110010";
                      t2addb <= "00110110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010110011";
                elsif cntr ="001010110011" THEN
                      t1addb <= "00110011";
                      t2addb <= "00110111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010110100";
                elsif cntr ="001010110100" THEN
                      t1addb <= "00110100";
                      t2addb <= "00110000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010110101";
                elsif cntr ="001010110101" THEN
                      t1addb <= "00110101";
                      t2addb <= "00110001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00101101";
                      cntr <= "001010110110";
                elsif cntr ="001010110110" THEN
                      t1addb <= "00110110";
                      t2addb <= "00110010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010110111";
                elsif cntr ="001010110111" THEN
                      t1addb <= "00110111";
                      t2addb <= "00110011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010111000";
                elsif cntr ="001010111000" THEN
                      t1addb <= "00111000";
                      t2addb <= "00111100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010111001";
                elsif cntr ="001010111001" THEN
                      t1addb <= "00111001";
                      t2addb <= "00111101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00101110";
                      cntr <= "001010111010";
                elsif cntr ="001010111010" THEN
                      t1addb <= "00111010";
                      t2addb <= "00111110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010111011";
                elsif cntr ="001010111011" THEN
                      t1addb <= "00111011";
                      t2addb <= "00111111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010111100";
                elsif cntr ="001010111100" THEN
                      t1addb <= "00111100";
                      t2addb <= "00111000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001010111101";
                elsif cntr ="001010111101" THEN
                      t1addb <= "00111101";
                      t2addb <= "00111001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00101111";
                      cntr <= "001010111110";
                elsif cntr ="001010111110" THEN
                      t1addb <= "00111110";
                      t2addb <= "00111010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001010111111";
                elsif cntr ="001010111111" THEN
                      t1addb <= "00111111";
                      t2addb <= "00111011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011000000";
                elsif cntr ="001011000000" THEN
                      t1addb <= "01000000";
                      t2addb <= "01000100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011000001";
                elsif cntr ="001011000001" THEN
                      t1addb <= "01000001";
                      t2addb <= "01000101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00110000";
                      cntr <= "001011000010";
                elsif cntr ="001011000010" THEN
                      t1addb <= "01000010";
                      t2addb <= "01000110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011000011";
                elsif cntr ="001011000011" THEN
                      t1addb <= "01000011";
                      t2addb <= "01000111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011000100";
                elsif cntr ="001011000100" THEN
                      t1addb <= "01000100";
                      t2addb <= "01000000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011000101";
                elsif cntr ="001011000101" THEN
                      t1addb <= "01000101";
                      t2addb <= "01000001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00110001";
                      cntr <= "001011000110";
                elsif cntr ="001011000110" THEN
                      t1addb <= "01000110";
                      t2addb <= "01000010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011000111";
                elsif cntr ="001011000111" THEN
                      t1addb <= "01000111";
                      t2addb <= "01000011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011001000";
                elsif cntr ="001011001000" THEN
                      t1addb <= "01001000";
                      t2addb <= "01001100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011001001";
                elsif cntr ="001011001001" THEN
                      t1addb <= "01001001";
                      t2addb <= "01001101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00110010";
                      cntr <= "001011001010";
                elsif cntr ="001011001010" THEN
                      t1addb <= "01001010";
                      t2addb <= "01001110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011001011";
                elsif cntr ="001011001011" THEN
                      t1addb <= "01001011";
                      t2addb <= "01001111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011001100";
                elsif cntr ="001011001100" THEN
                      t1addb <= "01001100";
                      t2addb <= "01001000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011001101";
                elsif cntr ="001011001101" THEN
                      t1addb <= "01001101";
                      t2addb <= "01001001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00110011";
                      cntr <= "001011001110";
                elsif cntr ="001011001110" THEN
                      t1addb <= "01001110";
                      t2addb <= "01001010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011001111";
                elsif cntr ="001011001111" THEN
                      t1addb <= "01001111";
                      t2addb <= "01001011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011010000";
                elsif cntr ="001011010000" THEN
                      t1addb <= "01010000";
                      t2addb <= "01010100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011010001";
                elsif cntr ="001011010001" THEN
                      t1addb <= "01010001";
                      t2addb <= "01010101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00110100";
                      cntr <= "001011010010";
                elsif cntr ="001011010010" THEN
                      t1addb <= "01010010";
                      t2addb <= "01010110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011010011";
                elsif cntr ="001011010011" THEN
                      t1addb <= "01010011";
                      t2addb <= "01010111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011010100";
                elsif cntr ="001011010100" THEN
                      t1addb <= "01010100";
                      t2addb <= "01010000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011010101";
                elsif cntr ="001011010101" THEN
                      t1addb <= "01010101";
                      t2addb <= "01010001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00110101";
                      cntr <= "001011010110";
                elsif cntr ="001011010110" THEN
                      t1addb <= "01010110";
                      t2addb <= "01010010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011010111";
                elsif cntr ="001011010111" THEN
                      t1addb <= "01010111";
                      t2addb <= "01010011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011011000";
                elsif cntr ="001011011000" THEN
                      t1addb <= "01011000";
                      t2addb <= "01011100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011011001";
                elsif cntr ="001011011001" THEN
                      t1addb <= "01011001";
                      t2addb <= "01011101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00110110";
                      cntr <= "001011011010";
                elsif cntr ="001011011010" THEN
                      t1addb <= "01011010";
                      t2addb <= "01011110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011011011";
                elsif cntr ="001011011011" THEN
                      t1addb <= "01011011";
                      t2addb <= "01011111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011011100";
                elsif cntr ="001011011100" THEN
                      t1addb <= "01011100";
                      t2addb <= "01011000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011011101";
                elsif cntr ="001011011101" THEN
                      t1addb <= "01011101";
                      t2addb <= "01011001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00110111";
                      cntr <= "001011011110";
                elsif cntr ="001011011110" THEN
                      t1addb <= "01011110";
                      t2addb <= "01011010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011011111";
                elsif cntr ="001011011111" THEN
                      t1addb <= "01011111";
                      t2addb <= "01011011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011100000";
                elsif cntr ="001011100000" THEN
                      t1addb <= "01100000";
                      t2addb <= "01100100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011100001";
                elsif cntr ="001011100001" THEN
                      t1addb <= "01100001";
                      t2addb <= "01100101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00111000";
                      cntr <= "001011100010";
                elsif cntr ="001011100010" THEN
                      t1addb <= "01100010";
                      t2addb <= "01100110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011100011";
                elsif cntr ="001011100011" THEN
                      t1addb <= "01100011";
                      t2addb <= "01100111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011100100";
                elsif cntr ="001011100100" THEN
                      t1addb <= "01100100";
                      t2addb <= "01100000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011100101";
                elsif cntr ="001011100101" THEN
                      t1addb <= "01100101";
                      t2addb <= "01100001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00111001";
                      cntr <= "001011100110";
                elsif cntr ="001011100110" THEN
                      t1addb <= "01100110";
                      t2addb <= "01100010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011100111";
                elsif cntr ="001011100111" THEN
                      t1addb <= "01100111";
                      t2addb <= "01100011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011101000";
                elsif cntr ="001011101000" THEN
                      t1addb <= "01101000";
                      t2addb <= "01101100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011101001";
                elsif cntr ="001011101001" THEN
                      t1addb <= "01101001";
                      t2addb <= "01101101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00111010";
                      cntr <= "001011101010";
                elsif cntr ="001011101010" THEN
                      t1addb <= "01101010";
                      t2addb <= "01101110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011101011";
                elsif cntr ="001011101011" THEN
                      t1addb <= "01101011";
                      t2addb <= "01101111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011101100";
                elsif cntr ="001011101100" THEN
                      t1addb <= "01101100";
                      t2addb <= "01101000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011101101";
                elsif cntr ="001011101101" THEN
                      t1addb <= "01101101";
                      t2addb <= "01101001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00111011";
                      cntr <= "001011101110";
                elsif cntr ="001011101110" THEN
                      t1addb <= "01101110";
                      t2addb <= "01101010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011101111";
                elsif cntr ="001011101111" THEN
                      t1addb <= "01101111";
                      t2addb <= "01101011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011110000";
                elsif cntr ="001011110000" THEN
                      t1addb <= "01110000";
                      t2addb <= "01110100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011110001";
                elsif cntr ="001011110001" THEN
                      t1addb <= "01110001";
                      t2addb <= "01110101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00111100";
                      cntr <= "001011110010";
                elsif cntr ="001011110010" THEN
                      t1addb <= "01110010";
                      t2addb <= "01110110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011110011";
                elsif cntr ="001011110011" THEN
                      t1addb <= "01110011";
                      t2addb <= "01110111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011110100";
                elsif cntr ="001011110100" THEN
                      t1addb <= "01110100";
                      t2addb <= "01110000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011110101";
                elsif cntr ="001011110101" THEN
                      t1addb <= "01110101";
                      t2addb <= "01110001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00111101";
                      cntr <= "001011110110";
                elsif cntr ="001011110110" THEN
                      t1addb <= "01110110";
                      t2addb <= "01110010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011110111";
                elsif cntr ="001011110111" THEN
                      t1addb <= "01110111";
                      t2addb <= "01110011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011111000";
                elsif cntr ="001011111000" THEN
                      t1addb <= "01111000";
                      t2addb <= "01111100";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011111001";
                elsif cntr ="001011111001" THEN
                      t1addb <= "01111001";
                      t2addb <= "01111101";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="00111110";
                      cntr <= "001011111010";
                elsif cntr ="001011111010" THEN
                      t1addb <= "01111010";
                      t2addb <= "01111110";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011111011";
                elsif cntr ="001011111011" THEN
                      t1addb <= "01111011";
                      t2addb <= "01111111";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011111100";
                elsif cntr ="001011111100" THEN
                      t1addb <= "01111100";
                      t2addb <= "01111000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      cntr <= "001011111101";
                elsif cntr ="001011111101" THEN
                      t1addb <= "01111101";
                      t2addb <= "01111001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="00111111";
                      cntr <= "001011111110";
                elsif cntr ="001011111110" THEN
                      t1addb <= "01111110";
                      t2addb <= "01111010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001011111111";
                elsif cntr ="001011111111" THEN
                      t1addb <= "01111111";
                      t2addb <= "01111011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      cntr <= "001100000000";
				elsif cntr ="001100000000" THEN
                      t1addb <= "10000000";
                      t2addb <= "10000010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                
                      
                      
                      
                      cntr <= "001100000001";
				elsif cntr ="001100000001" THEN
                      t1addb <= "10000001";
                      t2addb <= "10000011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                        zetain   <="01000000";      
                      cntr <= "001100000010";
                elsif cntr ="001100000010" THEN
                      t1addb <= "10000010";
                      t2addb <= "10000000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;      
                      
                      
                      
                            
                      cntr <= "001100000011";
                elsif cntr ="001100000011" THEN
                      t1addb <= "10000011";
                      t2addb <= "10000001";
                      bfrjin     <= t1doutb;      
                      bfrjplin <= t2doutb;      
                      
                      
                      
                        zetain   <="01000001";                  
                      cntr <= "001100000100";
                elsif cntr ="001100000100" THEN
                      t1addb <= "10000100";
                      t2addb <= "10000110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;      
                      
                      
                      
                                        
                      cntr <= "001100000101";
                elsif cntr ="001100000101" THEN
                      t1addb <= "10000101";
                      t2addb <= "10000111";
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      
                      
                      
                        zetain   <="01000010";                              
                      cntr <= "001100000110";   
                elsif cntr ="001100000110" THEN   
                      t1addb <= "10000110";
                      t2addb <= "10000100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;      
                      
                      
                      
                                                    
                      cntr <= "001100000111";  
                elsif cntr ="001100000111" THEN  
                      t1addb <= "10000111";
                      t2addb <= "10000101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                        zetain   <="01000011";                                         
                      cntr <= "001100001000";
                elsif cntr ="001100001000" THEN
                      t1addb <= "10001000";
                      t2addb <= "10001010";      
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      
                      
                      
                                                             
                      cntr <= "001100001001";
                elsif cntr ="001100001001" THEN
                      t1addb <= "10001001";
                      t2addb <= "10001011";
                      bfrjin     <= t2doutb;      
                      bfrjplin <= t1doutb;      
                      									
                
                
                      
                      
                        zetain   <="01000100";
                      cntr <= "001100001010";
                elsif cntr ="001100001010" THEN
                      t1addb <= "10001010";
                      t2addb <= "10001000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100001011";
                elsif cntr ="001100001011" THEN
                      t1addb <= "10001011";
                      t2addb <= "10001001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01000101";
                      cntr <= "001100001100";
                elsif cntr ="001100001100" THEN
                      t1addb <= "10001100";
                      t2addb <= "10001110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100001101";
                elsif cntr ="001100001101" THEN
                      t1addb <= "10001101";
                      t2addb <= "10001111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01000110";
                      cntr <= "001100001110";
                elsif cntr ="001100001110" THEN
                      t1addb <= "10001110";
                      t2addb <= "10001100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100001111";
                elsif cntr ="001100001111" THEN
                      t1addb <= "10001111";
                      t2addb <= "10001101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01000111";
                      cntr <= "001100010000";
                elsif cntr ="001100010000" THEN
                      t1addb <= "10010000";
                      t2addb <= "10010010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100010001";
                elsif cntr ="001100010001" THEN
                      t1addb <= "10010001";
                      t2addb <= "10010011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001000";
                      cntr <= "001100010010";
                elsif cntr ="001100010010" THEN
                      t1addb <= "10010010";
                      t2addb <= "10010000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100010011";
                elsif cntr ="001100010011" THEN
                      t1addb <= "10010011";
                      t2addb <= "10010001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001001";
                      cntr <= "001100010100";
                elsif cntr ="001100010100" THEN
                      t1addb <= "10010100";
                      t2addb <= "10010110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100010101";
                elsif cntr ="001100010101" THEN
                      t1addb <= "10010101";
                      t2addb <= "10010111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001010";
                      cntr <= "001100010110";
                elsif cntr ="001100010110" THEN
                      t1addb <= "10010110";
                      t2addb <= "10010100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100010111";
                elsif cntr ="001100010111" THEN
                      t1addb <= "10010111";
                      t2addb <= "10010101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001011";
                      cntr <= "001100011000";
                elsif cntr ="001100011000" THEN
                      t1addb <= "10011000";
                      t2addb <= "10011010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100011001";
                elsif cntr ="001100011001" THEN
                      t1addb <= "10011001";
                      t2addb <= "10011011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001100";
                      cntr <= "001100011010";
                elsif cntr ="001100011010" THEN
                      t1addb <= "10011010";
                      t2addb <= "10011000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100011011";
                elsif cntr ="001100011011" THEN
                      t1addb <= "10011011";
                      t2addb <= "10011001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001101";
                      cntr <= "001100011100";
                elsif cntr ="001100011100" THEN
                      t1addb <= "10011100";
                      t2addb <= "10011110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100011101";
                elsif cntr ="001100011101" THEN
                      t1addb <= "10011101";
                      t2addb <= "10011111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001110";
                      cntr <= "001100011110";
                elsif cntr ="001100011110" THEN
                      t1addb <= "10011110";
                      t2addb <= "10011100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100011111";
                elsif cntr ="001100011111" THEN
                      t1addb <= "10011111";
                      t2addb <= "10011101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01001111";
                      cntr <= "001100100000";
                elsif cntr ="001100100000" THEN
                      t1addb <= "10100000";
                      t2addb <= "10100010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100100001";
                elsif cntr ="001100100001" THEN
                      t1addb <= "10100001";
                      t2addb <= "10100011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010000";
                      cntr <= "001100100010";
                elsif cntr ="001100100010" THEN
                      t1addb <= "10100010";
                      t2addb <= "10100000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100100011";
                elsif cntr ="001100100011" THEN
                      t1addb <= "10100011";
                      t2addb <= "10100001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010001";
                      cntr <= "001100100100";
                elsif cntr ="001100100100" THEN
                      t1addb <= "10100100";
                      t2addb <= "10100110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100100101";
                elsif cntr ="001100100101" THEN
                      t1addb <= "10100101";
                      t2addb <= "10100111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010010";
                      cntr <= "001100100110";
                elsif cntr ="001100100110" THEN
                      t1addb <= "10100110";
                      t2addb <= "10100100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100100111";
                elsif cntr ="001100100111" THEN
                      t1addb <= "10100111";
                      t2addb <= "10100101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010011";
                      cntr <= "001100101000";
                elsif cntr ="001100101000" THEN
                      t1addb <= "10101000";
                      t2addb <= "10101010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100101001";
                elsif cntr ="001100101001" THEN
                      t1addb <= "10101001";
                      t2addb <= "10101011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010100";
                      cntr <= "001100101010";
                elsif cntr ="001100101010" THEN
                      t1addb <= "10101010";
                      t2addb <= "10101000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100101011";
                elsif cntr ="001100101011" THEN
                      t1addb <= "10101011";
                      t2addb <= "10101001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010101";
                      cntr <= "001100101100";
                elsif cntr ="001100101100" THEN
                      t1addb <= "10101100";
                      t2addb <= "10101110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100101101";
                elsif cntr ="001100101101" THEN
                      t1addb <= "10101101";
                      t2addb <= "10101111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010110";
                      cntr <= "001100101110";
                elsif cntr ="001100101110" THEN
                      t1addb <= "10101110";
                      t2addb <= "10101100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100101111";
                elsif cntr ="001100101111" THEN
                      t1addb <= "10101111";
                      t2addb <= "10101101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01010111";
                      cntr <= "001100110000";
                elsif cntr ="001100110000" THEN
                      t1addb <= "10110000";
                      t2addb <= "10110010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100110001";
                elsif cntr ="001100110001" THEN
                      t1addb <= "10110001";
                      t2addb <= "10110011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011000";
                      cntr <= "001100110010";
                elsif cntr ="001100110010" THEN
                      t1addb <= "10110010";
                      t2addb <= "10110000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100110011";
                elsif cntr ="001100110011" THEN
                      t1addb <= "10110011";
                      t2addb <= "10110001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011001";
                      cntr <= "001100110100";
                elsif cntr ="001100110100" THEN
                      t1addb <= "10110100";
                      t2addb <= "10110110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100110101";
                elsif cntr ="001100110101" THEN
                      t1addb <= "10110101";
                      t2addb <= "10110111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011010";
                      cntr <= "001100110110";
                elsif cntr ="001100110110" THEN
                      t1addb <= "10110110";
                      t2addb <= "10110100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100110111";
                elsif cntr ="001100110111" THEN
                      t1addb <= "10110111";
                      t2addb <= "10110101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011011";
                      cntr <= "001100111000";
                elsif cntr ="001100111000" THEN
                      t1addb <= "10111000";
                      t2addb <= "10111010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100111001";
                elsif cntr ="001100111001" THEN
                      t1addb <= "10111001";
                      t2addb <= "10111011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011100";
                      cntr <= "001100111010";
                elsif cntr ="001100111010" THEN
                      t1addb <= "10111010";
                      t2addb <= "10111000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100111011";
                elsif cntr ="001100111011" THEN
                      t1addb <= "10111011";
                      t2addb <= "10111001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011101";
                      cntr <= "001100111100";
                elsif cntr ="001100111100" THEN
                      t1addb <= "10111100";
                      t2addb <= "10111110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100111101";
                elsif cntr ="001100111101" THEN
                      t1addb <= "10111101";
                      t2addb <= "10111111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011110";
                      cntr <= "001100111110";
                elsif cntr ="001100111110" THEN
                      t1addb <= "10111110";
                      t2addb <= "10111100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001100111111";
                elsif cntr ="001100111111" THEN
                      t1addb <= "10111111";
                      t2addb <= "10111101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01011111";
                      cntr <= "001101000000";
                elsif cntr ="001101000000" THEN
                      t1addb <= "11000000";
                      t2addb <= "11000010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101000001";
                elsif cntr ="001101000001" THEN
                      t1addb <= "11000001";
                      t2addb <= "11000011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100000";
                      cntr <= "001101000010";
                elsif cntr ="001101000010" THEN
                      t1addb <= "11000010";
                      t2addb <= "11000000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101000011";
                elsif cntr ="001101000011" THEN
                      t1addb <= "11000011";
                      t2addb <= "11000001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100001";
                      cntr <= "001101000100";
                elsif cntr ="001101000100" THEN
                      t1addb <= "11000100";
                      t2addb <= "11000110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101000101";
                elsif cntr ="001101000101" THEN
                      t1addb <= "11000101";
                      t2addb <= "11000111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100010";
                      cntr <= "001101000110";
                elsif cntr ="001101000110" THEN
                      t1addb <= "11000110";
                      t2addb <= "11000100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101000111";
                elsif cntr ="001101000111" THEN
                      t1addb <= "11000111";
                      t2addb <= "11000101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100011";
                      cntr <= "001101001000";
                elsif cntr ="001101001000" THEN
                      t1addb <= "11001000";
                      t2addb <= "11001010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101001001";
                elsif cntr ="001101001001" THEN
                      t1addb <= "11001001";
                      t2addb <= "11001011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100100";
                      cntr <= "001101001010";
                elsif cntr ="001101001010" THEN
                      t1addb <= "11001010";
                      t2addb <= "11001000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101001011";
                elsif cntr ="001101001011" THEN
                      t1addb <= "11001011";
                      t2addb <= "11001001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100101";
                      cntr <= "001101001100";
                elsif cntr ="001101001100" THEN
                      t1addb <= "11001100";
                      t2addb <= "11001110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101001101";
                elsif cntr ="001101001101" THEN
                      t1addb <= "11001101";
                      t2addb <= "11001111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100110";
                      cntr <= "001101001110";
                elsif cntr ="001101001110" THEN
                      t1addb <= "11001110";
                      t2addb <= "11001100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101001111";
                elsif cntr ="001101001111" THEN
                      t1addb <= "11001111";
                      t2addb <= "11001101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01100111";
                      cntr <= "001101010000";
                elsif cntr ="001101010000" THEN
                      t1addb <= "11010000";
                      t2addb <= "11010010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101010001";
                elsif cntr ="001101010001" THEN
                      t1addb <= "11010001";
                      t2addb <= "11010011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101000";
                      cntr <= "001101010010";
                elsif cntr ="001101010010" THEN
                      t1addb <= "11010010";
                      t2addb <= "11010000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101010011";
                elsif cntr ="001101010011" THEN
                      t1addb <= "11010011";
                      t2addb <= "11010001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101001";
                      cntr <= "001101010100";
                elsif cntr ="001101010100" THEN
                      t1addb <= "11010100";
                      t2addb <= "11010110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101010101";
                elsif cntr ="001101010101" THEN
                      t1addb <= "11010101";
                      t2addb <= "11010111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101010";
                      cntr <= "001101010110";
                elsif cntr ="001101010110" THEN
                      t1addb <= "11010110";
                      t2addb <= "11010100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101010111";
                elsif cntr ="001101010111" THEN
                      t1addb <= "11010111";
                      t2addb <= "11010101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101011";
                      cntr <= "001101011000";
                elsif cntr ="001101011000" THEN
                      t1addb <= "11011000";
                      t2addb <= "11011010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101011001";
                elsif cntr ="001101011001" THEN
                      t1addb <= "11011001";
                      t2addb <= "11011011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101100";
                      cntr <= "001101011010";
                elsif cntr ="001101011010" THEN
                      t1addb <= "11011010";
                      t2addb <= "11011000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101011011";
                elsif cntr ="001101011011" THEN
                      t1addb <= "11011011";
                      t2addb <= "11011001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101101";
                      cntr <= "001101011100";
                elsif cntr ="001101011100" THEN
                      t1addb <= "11011100";
                      t2addb <= "11011110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101011101";
                elsif cntr ="001101011101" THEN
                      t1addb <= "11011101";
                      t2addb <= "11011111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101110";
                      cntr <= "001101011110";
                elsif cntr ="001101011110" THEN
                      t1addb <= "11011110";
                      t2addb <= "11011100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101011111";
                elsif cntr ="001101011111" THEN
                      t1addb <= "11011111";
                      t2addb <= "11011101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01101111";
                      cntr <= "001101100000";
                elsif cntr ="001101100000" THEN
                      t1addb <= "11100000";
                      t2addb <= "11100010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101100001";
                elsif cntr ="001101100001" THEN
                      t1addb <= "11100001";
                      t2addb <= "11100011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110000";
                      cntr <= "001101100010";
                elsif cntr ="001101100010" THEN
                      t1addb <= "11100010";
                      t2addb <= "11100000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101100011";
                elsif cntr ="001101100011" THEN
                      t1addb <= "11100011";
                      t2addb <= "11100001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110001";
                      cntr <= "001101100100";
                elsif cntr ="001101100100" THEN
                      t1addb <= "11100100";
                      t2addb <= "11100110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101100101";
                elsif cntr ="001101100101" THEN
                      t1addb <= "11100101";
                      t2addb <= "11100111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110010";
                      cntr <= "001101100110";
                elsif cntr ="001101100110" THEN
                      t1addb <= "11100110";
                      t2addb <= "11100100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101100111";
                elsif cntr ="001101100111" THEN
                      t1addb <= "11100111";
                      t2addb <= "11100101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110011";
                      cntr <= "001101101000";
                elsif cntr ="001101101000" THEN
                      t1addb <= "11101000";
                      t2addb <= "11101010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101101001";
                elsif cntr ="001101101001" THEN
                      t1addb <= "11101001";
                      t2addb <= "11101011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110100";
                      cntr <= "001101101010";
                elsif cntr ="001101101010" THEN
                      t1addb <= "11101010";
                      t2addb <= "11101000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101101011";
                elsif cntr ="001101101011" THEN
                      t1addb <= "11101011";
                      t2addb <= "11101001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110101";
                      cntr <= "001101101100";
                elsif cntr ="001101101100" THEN
                      t1addb <= "11101100";
                      t2addb <= "11101110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101101101";
                elsif cntr ="001101101101" THEN
                      t1addb <= "11101101";
                      t2addb <= "11101111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110110";
                      cntr <= "001101101110";
                elsif cntr ="001101101110" THEN
                      t1addb <= "11101110";
                      t2addb <= "11101100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101101111";
                elsif cntr ="001101101111" THEN
                      t1addb <= "11101111";
                      t2addb <= "11101101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01110111";
                      cntr <= "001101110000";
                elsif cntr ="001101110000" THEN
                      t1addb <= "11110000";
                      t2addb <= "11110010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101110001";
                elsif cntr ="001101110001" THEN
                      t1addb <= "11110001";
                      t2addb <= "11110011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111000";
                      cntr <= "001101110010";
                elsif cntr ="001101110010" THEN
                      t1addb <= "11110010";
                      t2addb <= "11110000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101110011";
                elsif cntr ="001101110011" THEN
                      t1addb <= "11110011";
                      t2addb <= "11110001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111001";
                      cntr <= "001101110100";
                elsif cntr ="001101110100" THEN
                      t1addb <= "11110100";
                      t2addb <= "11110110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101110101";
                elsif cntr ="001101110101" THEN
                      t1addb <= "11110101";
                      t2addb <= "11110111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111010";
                      cntr <= "001101110110";
                elsif cntr ="001101110110" THEN
                      t1addb <= "11110110";
                      t2addb <= "11110100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101110111";
                elsif cntr ="001101110111" THEN
                      t1addb <= "11110111";
                      t2addb <= "11110101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111011";
                      cntr <= "001101111000";
                elsif cntr ="001101111000" THEN
                      t1addb <= "11111000";
                      t2addb <= "11111010";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101111001";
                elsif cntr ="001101111001" THEN
                      t1addb <= "11111001";
                      t2addb <= "11111011";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111100";
                      cntr <= "001101111010";
                elsif cntr ="001101111010" THEN
                      t1addb <= "11111010";
                      t2addb <= "11111000";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101111011";
                elsif cntr ="001101111011" THEN
                      t1addb <= "11111011";
                      t2addb <= "11111001";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111101";
                      cntr <= "001101111100";
                elsif cntr ="001101111100" THEN
                      t1addb <= "11111100";
                      t2addb <= "11111110";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101111101";
                elsif cntr ="001101111101" THEN
                      t1addb <= "11111101";
                      t2addb <= "11111111";
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111110";
                      cntr <= "001101111110";
                elsif cntr ="001101111110" THEN
                      t1addb <= "11111110";
                      t2addb <= "11111100";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                      
                      cntr <= "001101111111";
                elsif cntr ="001101111111" THEN
                      t1addb <= "11111111";
                      t2addb <= "11111101";
                      bfrjin     <= t1doutb;
                      bfrjplin <= t2doutb;
                      
                      
                      
                      
                      
                        zetain   <="01111111";
                      cntr <= "001110000000";
                elsif cntr ="001110000000" THEN														
                      
                      
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                       
                      cntr <= "001110000001";
				elsif cntr ="001110000001" THEN						
                      
                      
                      bfrjin     <= t2doutb;
                      bfrjplin <= t1doutb;
                      
                      
                      
                      
                      
                       
                      cntr <= "001110000010";
                elsif cntr ="001110000010" THEN		      
                      
                      
                      
                      
                      
                      
                      
                            
                            
                             
                      cntr <= "001110000011";      
                elsif cntr ="001110000011" THEN		        
                      
                      
                      
                      
                      
                      
                      
                                  
                                  
                                   
                      cntr <= "001110000100";            
                elsif cntr ="001110000100" THEN		        
                      
                      
                      
                      
                      
                      
                      
                                        
                                        
                                         
                      cntr <= "001110000101";             
                elsif cntr ="001110000101" THEN		      
                      
                      
                      
                      
                      
                      
                      
                                               
                                               
                                                
                       cntr <= "001110000110";             
                 elsif cntr ="001110000110" THEN		      
                      
                      
                      
                      
                      
                      
                      
                                                     
                                                     
                                                      
                       cntr <= "001110000111";            
                 elsif cntr ="001110000111" THEN	      
                      
                      
                      
                      
                      
                      
                      
                                                           
                                                           
                                                           
                       cntr <= "001110001000";             
                 elsif cntr ="001110001000" THEN	       
                      
                      
                      
                      
                      
                      
                      
                                                           
                       
					
                                                           									
                       cntr <= "001110001001";       
                 elsif cntr ="001110001001" THEN	 

						
					  
					
				       cntr <= "001110001010";       
                 elsif cntr ="001110001010" THEN	 
					
					pdone <= '1';
					
					cntr <="001110001011";
				
				
				
				
				 elsif cntr ="001110001011" THEN	 

					cntr <="000000000000";
				
				
				END IF;
					
				
---------------------------------------------------------------------------------------------------------------------------------				
---------------------------------------------------------------------------------------------------------------------------------				
---------------------------------------------------------------------------------------------------------------------------------	

				
				
				
				IF cntr1 ="000000001001" THEN
					  	  					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00000000";
					  t2adda <= "00000000";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000001010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
					  t2adda <= "00000001";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000001011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
					  t2adda <= "00000010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000001100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
					  t2adda <= "00000011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000001101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00000100";
					  t2adda <= "00000100";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000001110" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
					  t2adda <= "00000101";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000001111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000010000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00000111";
					  t2adda <= "00000111";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000010001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00001000";
					  t2adda <= "00001000";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000010010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000010011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00001010";
					  t2adda <= "00001010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000010100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
					  t2adda <= "00001011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000010101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
					  t2adda <= "00001100";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000010110" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000010111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
					  t2adda <= "00001110";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000011000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00001111";
					  t2adda <= "00001111";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010000";
					  t2adda <= "00010000";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010001";
					  t2adda <= "00010001";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011011" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010010";
					  t2adda <= "00010010";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011100" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010011";
					  t2adda <= "00010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010100";
					  t2adda <= "00010100";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010101";
					  t2adda <= "00010101";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000011111" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010110";
					  t2adda <= "00010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000100000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00010111";
					  t2adda <= "00010111";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000100001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00011000";
					  t2adda <= "00011000";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000100010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000100011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000100100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
					  t2adda <= "00011011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000100101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00011100";
					  t2adda <= "00011100";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000100110" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00011101";
					  t2adda <= "00011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000100111" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00011110";
					  t2adda <= "00011110";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000101000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00011111";
					  t2adda <= "00011111";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000101001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00100000";
					  t2adda <= "00100000";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000101010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00100001";
					  t2adda <= "00100001";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000101011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000101100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
					  t2adda <= "00100011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000101101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000101110" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000101111" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00100110";
					  t2adda <= "00100110";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110000" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00100111";
					  t2adda <= "00100111";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000110010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00101001";
					  t2adda <= "00101001";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00101010";
					  t2adda <= "00101010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110100" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00101011";
					  t2adda <= "00101011";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00101100";
					  t2adda <= "00101100";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110110" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00101101";
					  t2adda <= "00101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000110111" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00101110";
					  t2adda <= "00101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000111000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00101111";
					  t2adda <= "00101111";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000111001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00110000";
					  t2adda <= "00110000";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000111010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00110001";
					  t2adda <= "00110001";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000000111011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
					  t2adda <= "00110010";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000111100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000000111101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
					  t2adda <= "00110100";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000111110" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
					  t2adda <= "00110101";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000000111111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
					  t2adda <= "00110110";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000001000000" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
					  
				elsif cntr1 ="000001000001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00111000";
					  t2adda <= "00111000";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001000010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
					  t2adda <= "00111001";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
					  
				      
				elsif cntr1 ="000001000011" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00111010";
					  t2adda <= "00111010";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001000100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "00111011";
					  t2adda <= "00111011";
					  t1dina <= bfrjout;
					  t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001000101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00111100";
					  t2adda <= "00111100";
					  t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001000110" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00111101";
					  t2adda <= "00111101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001000111" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00111110";
					  t2adda <= "00111110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001001000" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "00111111";
					  t2adda <= "00111111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000001001001" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000000";
					  t2adda <= "01000000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000001";
					  t2adda <= "01000001";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001011" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000010";
					  t2adda <= "01000010";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001100" THEN
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000011";
					  t2adda <= "01000011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000100";
					  t2adda <= "01000100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01000101";
					  t2adda <= "01000101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001001111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01000110";
					  t2adda <= "01000110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001010000" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
					  t2adda <= "01000111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001010001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01001000";
					  t2adda <= "01001000";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001010010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
					  t2adda <= "01001001";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001010011" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01001010";
					  t2adda <= "01001010";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001010100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
					  t2adda <= "01001011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001010101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01001100";
					  t2adda <= "01001100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001010110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01001101";
					  t2adda <= "01001101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001010111" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01001110";
					  t2adda <= "01001110";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001011000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01001111";
					  t2adda <= "01001111";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001011001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01010000";
					  t2adda <= "01010000";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001011010" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01010001";
					  t2adda <= "01010001";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001011011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
					  t2adda <= "01010010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001011100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010011";
					  t2adda <= "01010011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001011101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
					  t2adda <= "01010100";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001011110" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
					  t2adda <= "01010101";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001011111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
					  t2adda <= "01010110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100000" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
					  t2adda <= "01010111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
					  t2adda <= "01011000";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01011001";
					  t2adda <= "01011001";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001100011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
					  t2adda <= "01011010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
					  t2adda <= "01011011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
					  t2adda <= "01011100";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001100110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01011101";
					  t2adda <= "01011101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001100111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01011110";
					  t2adda <= "01011110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101000" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01011111";
					  t2adda <= "01011111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
					  t2adda <= "01100000";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001101010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
				elsif cntr1 ="000001101011" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01100010";
					  t2adda <= "01100010";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01100011";
					  t2adda <= "01100011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01100100";
					  t2adda <= "01100100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01100101";
					  t2adda <= "01100101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001101111" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01100110";
					  t2adda <= "01100110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001110000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01100111";
					  t2adda <= "01100111";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001110001" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
					  t2adda <= "01101000";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001110010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101001";
					  t2adda <= "01101001";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001110011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
					  t2adda <= "01101010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001110100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
					  t2adda <= "01101011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001110101" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
				elsif cntr1 ="000001110110" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01101101";
					  t2adda <= "01101101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001110111" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01101110";
					  t2adda <= "01101110";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111000" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01101111";
					  t2adda <= "01101111";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111001" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01110000";
					  t2adda <= "01110000";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111010" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01110001";
					  t2adda <= "01110001";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111011" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
					  t2adda <= "01110010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				elsif cntr1 ="000001111100" THEN
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01110011";
					  t2adda <= "01110011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111101" THEN
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01110100";
					  t2adda <= "01110100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111110" THEN
				      
					  
				
					  
					  
			
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01110101";
					  t2adda <= "01110101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000001111111" THEN
				      
					  
					  
					  
		
				      
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01110110";
					  t2adda <= "01110110";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000000" THEN
		
					  
				      
				      
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01110111";
					  t2adda <= "01110111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
				elsif cntr1 ="000010000001" THEN
				
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
				      t1adda <= "01111000";
				      t2adda <= "01111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000010" THEN

					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111001";
					  t2adda <= "01111001";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000011" THEN
					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111010";
					  t2adda <= "01111010";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000100" THEN

					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111011";
					  t2adda <= "01111011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000101" THEN
					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111100";
					  t2adda <= "01111100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000110" THEN

					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111101";
					  t2adda <= "01111101";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010000111" THEN

					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111110";
					  t2adda <= "01111110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010001000" THEN



					  
					  
					  
					  
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "01111111";
					  t2adda <= "01111111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				
				
				elsif cntr1 ="000010001001" THEN
					  t1wea <= '1';				
				      t2wea <= '1';
				      t1adda <= "10000000";
				      t2adda <= "10000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000001";
				      t2adda <= "10000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000010";
				      t2adda <= "10000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000011";
				      t2adda <= "10000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000100";
				      t2adda <= "10000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000101";
				      t2adda <= "10000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010001111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000110";
				      t2adda <= "10000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000111";
				      t2adda <= "10000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001000";
				      t2adda <= "10001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001001";
				      t2adda <= "10001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001010";
				      t2adda <= "10001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001011";
				      t2adda <= "10001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001100";
				      t2adda <= "10001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001101";
				      t2adda <= "10001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010010111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001110";
				      t2adda <= "10001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001111";
				      t2adda <= "10001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010000";
				      t2adda <= "10010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010001";
				      t2adda <= "10010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010010";
				      t2adda <= "10010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010011";
				      t2adda <= "10010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010100";
				      t2adda <= "10010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010101";
				      t2adda <= "10010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010011111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010110";
				      t2adda <= "10010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010111";
				      t2adda <= "10010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011000";
				      t2adda <= "10011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011001";
				      t2adda <= "10011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011010";
				      t2adda <= "10011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011011";
				      t2adda <= "10011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011100";
				      t2adda <= "10011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011101";
				      t2adda <= "10011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010100111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011110";
				      t2adda <= "10011110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011111";
				      t2adda <= "10011111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100000";
				      t2adda <= "10100000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100001";
				      t2adda <= "10100001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100010";
				      t2adda <= "10100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100011";
				      t2adda <= "10100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100100";
				      t2adda <= "10100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100101";
				      t2adda <= "10100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010101111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100110";
				      t2adda <= "10100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100111";
				      t2adda <= "10100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101000";
				      t2adda <= "10101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101001";
				      t2adda <= "10101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101010";
				      t2adda <= "10101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101011";
				      t2adda <= "10101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101100";
				      t2adda <= "10101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101101";
				      t2adda <= "10101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010110111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101110";
				      t2adda <= "10101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101111";
				      t2adda <= "10101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110000";
				      t2adda <= "10110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110001";
				      t2adda <= "10110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110010";
				      t2adda <= "10110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110011";
				      t2adda <= "10110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110100";
				      t2adda <= "10110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110101";
				      t2adda <= "10110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000010111111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110110";
				      t2adda <= "10110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
					  
				elsif cntr1 ="000011000000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110111";
				      t2adda <= "10110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011000001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111000";
				      t2adda <= "10111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				elsif cntr1 ="000011000010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111001";
				      t2adda <= "10111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
					  
					  
				elsif cntr1 ="000011000011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111010";
				      t2adda <= "10111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011000100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111011";
				      t2adda <= "10111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011000101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111100";
				      t2adda <= "10111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011000110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111101";
				      t2adda <= "10111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011000111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111110";
				      t2adda <= "10111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111111";
				      t2adda <= "10111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000000";
				      t2adda <= "11000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000001";
				      t2adda <= "11000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000010";
				      t2adda <= "11000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000011";
				      t2adda <= "11000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000100";
				      t2adda <= "11000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000101";
				      t2adda <= "11000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011001111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000110";
				      t2adda <= "11000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000111";
				      t2adda <= "11000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001000";
				      t2adda <= "11001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001001";
				      t2adda <= "11001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001010";
				      t2adda <= "11001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001011";
				      t2adda <= "11001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001100";
				      t2adda <= "11001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001101";
				      t2adda <= "11001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011010111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001110";
				      t2adda <= "11001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001111";
				      t2adda <= "11001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010000";
				      t2adda <= "11010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010001";
				      t2adda <= "11010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010010";
				      t2adda <= "11010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010011";
				      t2adda <= "11010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010100";
				      t2adda <= "11010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010101";
				      t2adda <= "11010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011011111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010110";
				      t2adda <= "11010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010111";
				      t2adda <= "11010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011000";
				      t2adda <= "11011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011001";
				      t2adda <= "11011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011010";
				      t2adda <= "11011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011011";
				      t2adda <= "11011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011100";
				      t2adda <= "11011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011101";
				      t2adda <= "11011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011100111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011110";
				      t2adda <= "11011110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011111";
				      t2adda <= "11011111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100000";
				      t2adda <= "11100000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
			          
				elsif cntr1 ="000011101010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100001";
				      t2adda <= "11100001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101011" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100010";
				      t2adda <= "11100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101100" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100011";
				      t2adda <= "11100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101101" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100100";
				      t2adda <= "11100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101110" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100101";
				      t2adda <= "11100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011101111" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100110";
				      t2adda <= "11100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011110000" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100111";
				      t2adda <= "11100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011110001" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101000";
				      t2adda <= "11101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011110010" THEN
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101001";
				      t2adda <= "11101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				      
				      
				elsif cntr1 ="000011110011" THEN
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101010";
					  t2adda <= "11101010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
					  
					  
					  
				elsif cntr1 ="000011110100" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11101011";
				      t2adda <= "11101011";
				      t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
					  
					  
					  
				elsif cntr1 ="000011110101" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11101100";
					  t2adda <= "11101100";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
					  
					  
					  
					  
				elsif cntr1 ="000011110110" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11101101";
					  t2adda <= "11101101";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
				      
				      
					  
					  
				elsif cntr1 ="000011110111" THEN
				      t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11101110";
					  t2adda <= "11101110";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
					  
				      
				      
				elsif cntr1 ="000011111000" THEN
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101111";
					  t2adda <= "11101111";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
					  
					  
					  
				elsif cntr1 ="000011111001" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11110000";
				      t2adda <= "11110000";
				      t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  
					  
					  
					  
					  
				elsif cntr1 ="000011111010" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11110001";
					  t2adda <= "11110001";
					  t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
					  
					  
					  
					  
				elsif cntr1 ="000011111011" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11110010";
					  t2adda <= "11110010";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
					  	
					  
					  
					  
					  
				elsif cntr1 ="000011111100" THEN
					  t1wea <= '1';
					  t2wea <= '1';
					  t1adda <= "11110011";
					  t2adda <= "11110011";
					  t1dina <= bfrjplout;
					  t2dina <= bfrjout;
				      
                      
                      
                      
                      
                elsif cntr1 ="000011111101" THEN
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110100";
                      t2adda <= "11110100";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                      
                      
                elsif cntr1 ="000011111110" THEN
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110101";
                      t2adda <= "11110101";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                      
                elsif cntr1 ="000011111111" THEN
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110110";
                      t2adda <= "11110110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
				elsif cntr1 ="000100000000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110111";
                      t2adda <= "11110111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
			          
                
                elsif cntr1 ="000100000001" THEN
                
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111000";
                      t2adda <= "11111000";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
				      
				elsif cntr1 ="000100000010" THEN
                      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111001";
				      t2adda <= "11111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				             
				            
                
                elsif cntr1 ="000100000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111010";
				      t2adda <= "11111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                   
				                  
				
				elsif cntr1 ="000100000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111011";
				      t2adda <= "11111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                         
				                        
				
				elsif cntr1 ="000100000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111100";
				      t2adda <= "11111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                               
				                              
				
				elsif cntr1 ="000100000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111101";
				      t2adda <= "11111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                     
				                                    
				
				elsif cntr1 ="000100000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111110";
				      t2adda <= "11111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                       
				                                       
				
				elsif cntr1 ="000100001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111111";
				      t2adda <= "11111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                   
				                                   
				
				elsif cntr1 ="000100001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000000";
				      t2adda <= "00000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
				      t2adda <= "00000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001011" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
				      t2adda <= "00000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
				      t2adda <= "00000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000100";
				      t2adda <= "00000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
				      t2adda <= "00000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000111";
				      t2adda <= "00000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="000100010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001000";
				      t2adda <= "00001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
                      
				elsif cntr1 ="000100010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001010";
				      t2adda <= "00001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
				      t2adda <= "00001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000100010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
				      t2adda <= "00001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
				      t2adda <= "00001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "00001111";
				      t2adda <= "00001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010000";
				      t2adda <= "00010000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011010" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010001";
				      t2adda <= "00010001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010010";
				      t2adda <= "00010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011100" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010011";
				      t2adda <= "00010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010100";
				      t2adda <= "00010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010101";
				      t2adda <= "00010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010110";
				      t2adda <= "00010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010111";
				      t2adda <= "00010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011000";
				      t2adda <= "00011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                elsif cntr1 ="000100100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000100100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
				      t2adda <= "00011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011100";
				      t2adda <= "00011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000100100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011101";
				      t2adda <= "00011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011110";
				      t2adda <= "00011110";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011111";
				      t2adda <= "00011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "00100000";
				      t2adda <= "00100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100001";
				      t2adda <= "00100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101011" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
				      t2adda <= "00100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101101" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100110";
				      t2adda <= "00100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100111";
				      t2adda <= "00100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101001";
				      t2adda <= "00101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="000100110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101010";
				      t2adda <= "00101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101011";
				      t2adda <= "00101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
                      
				elsif cntr1 ="000100110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101100";
				      t2adda <= "00101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101101";
				      t2adda <= "00101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000100110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101110";
				      t2adda <= "00101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101111";
				      t2adda <= "00101111";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110000";
				      t2adda <= "00110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "00110001";
				      t2adda <= "00110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
				      t2adda <= "00110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111100" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
				      t2adda <= "00110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111110" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
				      t2adda <= "00110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
				      t2adda <= "00110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111000";
				      t2adda <= "00111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
				      t2adda <= "00111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111010";
				      t2adda <= "00111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="000101000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111011";
				      t2adda <= "00111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111100";
				      t2adda <= "00111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000101000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111101";
				      t2adda <= "00111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111110";
				      t2adda <= "00111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000101001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111111";
				      t2adda <= "00111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000000";
				      t2adda <= "01000000";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000001";
				      t2adda <= "01000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "01000010";
				      t2adda <= "01000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000011";
				      t2adda <= "01000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001101" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000100";
				      t2adda <= "01000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000101";
				      t2adda <= "01000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001111" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000110";
				      t2adda <= "01000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
				      t2adda <= "01000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001000";
				      t2adda <= "01001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
				      t2adda <= "01001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001010";
				      t2adda <= "01001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
				      t2adda <= "01001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="000101010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001100";
				      t2adda <= "01001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001101";
				      t2adda <= "01001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
                      
				elsif cntr1 ="000101010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001110";
				      t2adda <= "01001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001111";
				      t2adda <= "01001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000101011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010000";
				      t2adda <= "01010000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010001";
				      t2adda <= "01010001";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
				      t2adda <= "01010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "01010011";
				      t2adda <= "01010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
				      t2adda <= "01010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011110" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
				      t2adda <= "01010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
				      t2adda <= "01010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100000" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
				      t2adda <= "01010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
				      t2adda <= "01011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011001";
				      t2adda <= "01011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
				      t2adda <= "01011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
				      t2adda <= "01011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
				      t2adda <= "01011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="000101100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011101";
				      t2adda <= "01011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011110";
				      t2adda <= "01011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000101101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011111";
				      t2adda <= "01011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
				      t2adda <= "01100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000101101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100010";
				      t2adda <= "01100010";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100011";
				      t2adda <= "01100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "01100100";
				      t2adda <= "01100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100101";
				      t2adda <= "01100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101111" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100110";
				      t2adda <= "01100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100111";
				      t2adda <= "01100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110001" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
				      t2adda <= "01101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101001";
				      t2adda <= "01101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
				      t2adda <= "01101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
				      t2adda <= "01101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101101";
				      t2adda <= "01101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="000101110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101110";
				      t2adda <= "01101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101111";
				      t2adda <= "01101111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
                      
				elsif cntr1 ="000101111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110000";
				      t2adda <= "01110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110001";
				      t2adda <= "01110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000101111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
				      t2adda <= "01110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110011";
				      t2adda <= "01110011";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110100";
				      t2adda <= "01110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "01110101";
				      t2adda <= "01110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110110";
				      t2adda <= "01110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110111";
				      t2adda <= "01110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110000001" THEN
				
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111000";
				      t2adda <= "01111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110000010" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111001";
				      t2adda <= "01111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="000110000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111010";
				      t2adda <= "01111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
                
                elsif cntr1 ="000110000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111011";
				      t2adda <= "01111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				
				elsif cntr1 ="000110000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111100";
				      t2adda <= "01111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				
				elsif cntr1 ="000110000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111101";
				      t2adda <= "01111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				
				elsif cntr1 ="000110000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111110";
				      t2adda <= "01111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                        
				                                        
				  
				elsif cntr1 ="000110001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111111";
				      t2adda <= "01111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                
				                                
				
				elsif cntr1 ="000110001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000000";
				      t2adda <= "10000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000001";
				      t2adda <= "10000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000010";
				      t2adda <= "10000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				      
				elsif cntr1 ="000110001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000011";
				      t2adda <= "10000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001101" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "10000100";
				      t2adda <= "10000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000101";
				      t2adda <= "10000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000110";
				      t2adda <= "10000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000111";
				      t2adda <= "10000111";
				      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001000";
				      t2adda <= "10001000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110010010" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001001";
				      t2adda <= "10001001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001010";
				      t2adda <= "10001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001011";
				      t2adda <= "10001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "10001100";
				      t2adda <= "10001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001101";
				      t2adda <= "10001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001110";
				      t2adda <= "10001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001111";
				      t2adda <= "10001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000110011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010000";
				      t2adda <= "10010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011010" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010001";
				      t2adda <= "10010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010010";
				      t2adda <= "10010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="000110011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010011";
				      t2adda <= "10010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010100";
                      t2adda <= "10010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010101";
				      t2adda <= "10010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010110";
				      t2adda <= "10010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010111";
				      t2adda <= "10010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				      
				elsif cntr1 ="000110100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011000";
				      t2adda <= "10011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110100010" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011001";
				      t2adda <= "10011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011010";
				      t2adda <= "10011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011011";
				      t2adda <= "10011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011100";
				      t2adda <= "10011100";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011101";
				      t2adda <= "10011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011110";
				      t2adda <= "10011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011111";
				      t2adda <= "10011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000110101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100000";
				      t2adda <= "10100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101010" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "10100001";
				      t2adda <= "10100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100010";
				      t2adda <= "10100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100011";
				      t2adda <= "10100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100100";
				      t2adda <= "10100100";
				      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100101";
				      t2adda <= "10100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101111" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100110";
				      t2adda <= "10100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100111";
				      t2adda <= "10100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101000";
				      t2adda <= "10101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "10101001";
				      t2adda <= "10101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101010";
				      t2adda <= "10101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101011";
				      t2adda <= "10101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101100";
				      t2adda <= "10101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000110110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101101";
				      t2adda <= "10101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110110111" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101110";
				      t2adda <= "10101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101111";
				      t2adda <= "10101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="000110111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110000";
				      t2adda <= "10110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110001";
                      t2adda <= "10110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110010";
				      t2adda <= "10110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110011";
				      t2adda <= "10110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110100";
				      t2adda <= "10110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				      
				elsif cntr1 ="000110111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110101";
				      t2adda <= "10110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111111" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110110";
				      t2adda <= "10110110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110111";
				      t2adda <= "10110111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111000";
				      t2adda <= "10111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111001";
				      t2adda <= "10111001";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111010";
				      t2adda <= "10111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111011";
				      t2adda <= "10111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111100";
				      t2adda <= "10111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000111000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111101";
				      t2adda <= "10111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000111" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "10111110";
				      t2adda <= "10111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111111";
				      t2adda <= "10111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000000";
				      t2adda <= "11000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000001";
				      t2adda <= "11000001";
				      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000010";
				      t2adda <= "11000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001100" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000011";
				      t2adda <= "11000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000100";
				      t2adda <= "11000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000101";
				      t2adda <= "11000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "11000110";
				      t2adda <= "11000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000111";
				      t2adda <= "11000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001000";
				      t2adda <= "11001000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001001";
				      t2adda <= "11001001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                      
				      
				      
				elsif cntr1 ="000111010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001010";
				      t2adda <= "11001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111010100" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001011";
				      t2adda <= "11001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001100";
				      t2adda <= "11001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="000111010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001101";
				      t2adda <= "11001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001110";
                      t2adda <= "11001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001111";
				      t2adda <= "11001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010000";
				      t2adda <= "11010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010001";
				      t2adda <= "11010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				      
				elsif cntr1 ="000111011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010010";
				      t2adda <= "11010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011100" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010011";
				      t2adda <= "11010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010100";
				      t2adda <= "11010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010101";
				      t2adda <= "11010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010110";
				      t2adda <= "11010110";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010111";
				      t2adda <= "11010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011000";
				      t2adda <= "11011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011001";
				      t2adda <= "11011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="000111100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011010";
				      t2adda <= "11011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100100" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "11011011";
				      t2adda <= "11011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011100";
				      t2adda <= "11011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011101";
				      t2adda <= "11011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011110";
				      t2adda <= "11011110";
				      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011111";
				      t2adda <= "11011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111101001" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100000";
				      t2adda <= "11100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100001";
				      t2adda <= "11100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100010";
				      t2adda <= "11100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100011";
				      t2adda <= "11100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000111101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100100";
				      t2adda <= "11100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100101";
				      t2adda <= "11100101";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100110";
				      t2adda <= "11100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "11100111";
				      t2adda <= "11100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101000";
				      t2adda <= "11101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111110010" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101001";
				      t2adda <= "11101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101010";
				      t2adda <= "11101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111110100" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101011";
				      t2adda <= "11101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101100";
				      t2adda <= "11101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101101";
				      t2adda <= "11101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101110";
				      t2adda <= "11101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101111";
                      t2adda <= "11101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110000";
				      t2adda <= "11110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111010" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "11110001";
				      t2adda <= "11110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110010";
				      t2adda <= "11110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111100" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110011";
				      t2adda <= "11110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110100";
				      t2adda <= "11110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110101";
				      t2adda <= "11110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="000111111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110110";
				      t2adda <= "11110110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110111";
				      t2adda <= "11110111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111000";
                      t2adda <= "11111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="001000000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111001";
				      t2adda <= "11111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="001000000011" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "11111010";
				      t2adda <= "11111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				elsif cntr1 ="001000000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111011";
				      t2adda <= "11111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				elsif cntr1 ="001000000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111100";
				      t2adda <= "11111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
                                              
				elsif cntr1 ="001000000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111101";
				      t2adda <= "11111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				
				elsif cntr1 ="001000000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111110";
				      t2adda <= "11111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
                                                          
				                                          
				    
				elsif cntr1 ="001000001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111111";
				      t2adda <= "11111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                 
				                                 
				
				elsif cntr1 ="001000001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000000";
				      t2adda <= "00000000";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
				      t2adda <= "00000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
				      t2adda <= "00000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
				      t2adda <= "00000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000100";
				      t2adda <= "00000100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
				      t2adda <= "00000101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
                      
				      
				elsif cntr1 ="001000010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000111";
				      t2adda <= "00000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001000";
				      t2adda <= "00001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001010";
				      t2adda <= "00001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
				      t2adda <= "00001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
				      t2adda <= "00001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="001000010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
				      t2adda <= "00001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000011000" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001111";
				      t2adda <= "00001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010000";
				      t2adda <= "00010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010001";
				      t2adda <= "00010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010010";
				      t2adda <= "00010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010011";
				      t2adda <= "00010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010100";
				      t2adda <= "00010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "00010101";
				      t2adda <= "00010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010110";
				      t2adda <= "00010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000100000" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010111";
				      t2adda <= "00010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011000";
				      t2adda <= "00011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000100010" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
				      t2adda <= "00011011";
				      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011100";
				      t2adda <= "00011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011101";
                      t2adda <= "00011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011110";
				      t2adda <= "00011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101000" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "00011111";
				      t2adda <= "00011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100000";
				      t2adda <= "00100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100001";
				      t2adda <= "00100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
                      
				elsif cntr1 ="001000101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
				      t2adda <= "00100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				      
				elsif cntr1 ="001000101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
                      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100110";
				      t2adda <= "00100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100111";
				      t2adda <= "00100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101001";
				      t2adda <= "00101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101010";
				      t2adda <= "00101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101011";
				      t2adda <= "00101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				      
				elsif cntr1 ="001000110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101100";
				      t2adda <= "00101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101101";
				      t2adda <= "00101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101110";
				      t2adda <= "00101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101111";
				      t2adda <= "00101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110000";
				      t2adda <= "00110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110001";
				      t2adda <= "00110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
                elsif cntr1 ="001000111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
				      t2adda <= "00110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111101" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
				      t2adda <= "00110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
				      t2adda <= "00110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
				      t2adda <= "00110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111000";
				      t2adda <= "00111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
				      t2adda <= "00111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "00111010";
				      t2adda <= "00111010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111011";
				      t2adda <= "00111011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000101" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111100";
				      t2adda <= "00111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111101";
				      t2adda <= "00111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000111" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111110";
				      t2adda <= "00111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111111";
				      t2adda <= "00111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000000";
				      t2adda <= "01000000";
				      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000001";
				      t2adda <= "01000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000010";
                      t2adda <= "01000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000011";
				      t2adda <= "01000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001101" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "01000100";
				      t2adda <= "01000100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000101";
				      t2adda <= "01000101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000110";
				      t2adda <= "01000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
                      
				elsif cntr1 ="001001010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
				      t2adda <= "01000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001000";
				      t2adda <= "01001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
                      
				      
				elsif cntr1 ="001001010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
				      t2adda <= "01001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001010";
				      t2adda <= "01001010";
                      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
				      t2adda <= "01001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001100";
				      t2adda <= "01001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001101";
				      t2adda <= "01001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001110";
				      t2adda <= "01001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001111";
				      t2adda <= "01001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010000";
				      t2adda <= "01010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
                      
				elsif cntr1 ="001001011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010001";
				      t2adda <= "01010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
				      t2adda <= "01010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010011";
				      t2adda <= "01010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
				      t2adda <= "01010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
				      t2adda <= "01010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
				      t2adda <= "01010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
                elsif cntr1 ="001001100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
				      t2adda <= "01010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
				      t2adda <= "01011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001100010" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011001";
				      t2adda <= "01011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
				      t2adda <= "01011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
				      t2adda <= "01011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
				      t2adda <= "01011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011101";
				      t2adda <= "01011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011110";
				      t2adda <= "01011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
                      t1adda <= "01011111";
				      t2adda <= "01011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
				      t2adda <= "01100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001101010" THEN
				      
				      
                      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100010";
				      t2adda <= "01100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101100" THEN
                      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100011";
				      t2adda <= "01100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100100";
				      t2adda <= "01100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100101";
				      t2adda <= "01100101";
				      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100110";
				      t2adda <= "01100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100111";
                      t2adda <= "01100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
				      t2adda <= "01101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001110010" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
				      t1adda <= "01101001";
				      t2adda <= "01101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
				      t2adda <= "01101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110100" THEN
				      
                      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
				      t2adda <= "01101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101101";
				      t2adda <= "01101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101110";
				      t2adda <= "01101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101111";
				      t2adda <= "01101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110000";
				      t2adda <= "01110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110001";
				      t2adda <= "01110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
				      t2adda <= "01110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110011";
				      t2adda <= "01110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110100";
				      t2adda <= "01110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
                      
				      
				elsif cntr1 ="001001111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110101";
				      t2adda <= "01110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110110";
				      t2adda <= "01110110";
				      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110111";
				      t2adda <= "01110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111000";
                      t2adda <= "01111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001010000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111001";
				      t2adda <= "01111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				            
				            
				
				elsif cntr1 ="001010000011" THEN
				      
				      
				      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111010";
                      t2adda <= "01111010";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                                  
                                  
                                  
                elsif cntr1 ="001010000100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111011";
                      t2adda <= "01111011";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                                        
                                        
                
                elsif cntr1 ="001010000101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111100";
                      t2adda <= "01111100";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                              
                                              
                elsif cntr1 ="001010000110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111101";
                      t2adda <= "01111101";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                                    
                                                    
                
                elsif cntr1 ="001010000111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111110";
                      t2adda <= "01111110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                                       
                                                       
                
                elsif cntr1 ="001010001000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "01111111";
                      t2adda <= "01111111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                                       
                                                       
                
                elsif cntr1 ="001010001001" THEN				
                
                
					  t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000000";
                      t2adda <= "10000000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010001010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000001";
                      t2adda <= "10000001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010001011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000010";
                      t2adda <= "10000010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010001100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000011";
                      t2adda <= "10000011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010001101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000100";
                      t2adda <= "10000100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010001110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000101";
                      t2adda <= "10000101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010001111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000110";
                      t2adda <= "10000110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010010000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10000111";
                      t2adda <= "10000111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010010001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001000";
                      t2adda <= "10001000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010010010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001001";
                      t2adda <= "10001001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010010011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001010";
                      t2adda <= "10001010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010010100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001011";
                      t2adda <= "10001011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010010101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001100";
                      t2adda <= "10001100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010010110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001101";
                      t2adda <= "10001101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010010111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001110";
                      t2adda <= "10001110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010011000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10001111";
                      t2adda <= "10001111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010011001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010000";
                      t2adda <= "10010000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010011010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010001";
                      t2adda <= "10010001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010011011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010010";
                      t2adda <= "10010010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010011100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010011";
                      t2adda <= "10010011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010011101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010100";
                      t2adda <= "10010100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010011110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010101";
                      t2adda <= "10010101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010011111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010110";
                      t2adda <= "10010110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010100000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10010111";
                      t2adda <= "10010111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010100001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011000";
                      t2adda <= "10011000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010100010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011001";
                      t2adda <= "10011001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010100011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011010";
                      t2adda <= "10011010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010100100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011011";
                      t2adda <= "10011011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010100101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011100";
                      t2adda <= "10011100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010100110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011101";
                      t2adda <= "10011101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010100111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011110";
                      t2adda <= "10011110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010101000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10011111";
                      t2adda <= "10011111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010101001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100000";
                      t2adda <= "10100000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010101010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100001";
                      t2adda <= "10100001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010101011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100010";
                      t2adda <= "10100010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010101100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100011";
                      t2adda <= "10100011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010101101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100100";
                      t2adda <= "10100100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010101110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100101";
                      t2adda <= "10100101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010101111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100110";
                      t2adda <= "10100110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010110000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10100111";
                      t2adda <= "10100111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010110001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101000";
                      t2adda <= "10101000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010110010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101001";
                      t2adda <= "10101001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010110011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101010";
                      t2adda <= "10101010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010110100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101011";
                      t2adda <= "10101011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010110101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101100";
                      t2adda <= "10101100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010110110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101101";
                      t2adda <= "10101101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010110111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101110";
                      t2adda <= "10101110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010111000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10101111";
                      t2adda <= "10101111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010111001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110000";
                      t2adda <= "10110000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010111010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110001";
                      t2adda <= "10110001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010111011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110010";
                      t2adda <= "10110010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010111100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110011";
                      t2adda <= "10110011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001010111101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110100";
                      t2adda <= "10110100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001010111110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110101";
                      t2adda <= "10110101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001010111111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110110";
                      t2adda <= "10110110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011000000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10110111";
                      t2adda <= "10110111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011000001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111000";
                      t2adda <= "10111000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011000010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111001";
                      t2adda <= "10111001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011000011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111010";
                      t2adda <= "10111010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011000100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111011";
                      t2adda <= "10111011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011000101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111100";
                      t2adda <= "10111100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011000110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111101";
                      t2adda <= "10111101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011000111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111110";
                      t2adda <= "10111110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011001000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "10111111";
                      t2adda <= "10111111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011001001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000000";
                      t2adda <= "11000000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011001010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000001";
                      t2adda <= "11000001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011001011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000010";
                      t2adda <= "11000010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011001100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000011";
                      t2adda <= "11000011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011001101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000100";
                      t2adda <= "11000100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011001110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000101";
                      t2adda <= "11000101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011001111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000110";
                      t2adda <= "11000110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011010000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11000111";
                      t2adda <= "11000111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011010001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001000";
                      t2adda <= "11001000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011010010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001001";
                      t2adda <= "11001001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011010011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001010";
                      t2adda <= "11001010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011010100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001011";
                      t2adda <= "11001011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011010101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001100";
                      t2adda <= "11001100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011010110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001101";
                      t2adda <= "11001101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011010111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001110";
                      t2adda <= "11001110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011011000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11001111";
                      t2adda <= "11001111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011011001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010000";
                      t2adda <= "11010000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011011010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010001";
                      t2adda <= "11010001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011011011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010010";
                      t2adda <= "11010010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011011100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010011";
                      t2adda <= "11010011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011011101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010100";
                      t2adda <= "11010100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011011110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010101";
                      t2adda <= "11010101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011011111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010110";
                      t2adda <= "11010110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011100000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11010111";
                      t2adda <= "11010111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011100001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011000";
                      t2adda <= "11011000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011100010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011001";
                      t2adda <= "11011001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011100011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011010";
                      t2adda <= "11011010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011100100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011011";
                      t2adda <= "11011011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011100101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011100";
                      t2adda <= "11011100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011100110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011101";
                      t2adda <= "11011101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011100111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011110";
                      t2adda <= "11011110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011101000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11011111";
                      t2adda <= "11011111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011101001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100000";
                      t2adda <= "11100000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011101010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100001";
                      t2adda <= "11100001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011101011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100010";
                      t2adda <= "11100010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011101100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100011";
                      t2adda <= "11100011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011101101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100100";
                      t2adda <= "11100100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011101110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100101";
                      t2adda <= "11100101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011101111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100110";
                      t2adda <= "11100110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011110000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11100111";
                      t2adda <= "11100111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011110001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101000";
                      t2adda <= "11101000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011110010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101001";
                      t2adda <= "11101001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011110011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101010";
                      t2adda <= "11101010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011110100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101011";
                      t2adda <= "11101011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011110101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101100";
                      t2adda <= "11101100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011110110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101101";
                      t2adda <= "11101101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011110111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101110";
                      t2adda <= "11101110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011111000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11101111";
                      t2adda <= "11101111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011111001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110000";
                      t2adda <= "11110000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011111010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110001";
                      t2adda <= "11110001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011111011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110010";
                      t2adda <= "11110010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011111100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110011";
                      t2adda <= "11110011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
                elsif cntr1 ="001011111101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110100";
                      t2adda <= "11110100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001011111110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110101";
                      t2adda <= "11110101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001011111111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110110";
                      t2adda <= "11110110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
				elsif cntr1 ="001100000000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11110111";
                      t2adda <= "11110111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                      
                      
                      
				elsif cntr1 ="001100000001" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111000";
                      t2adda <= "11111000";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                      
                      
                elsif cntr1 ="001100000010" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111001";
                      t2adda <= "11111001";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                            
                            
                            
                elsif cntr1 ="001100000011" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111010";
                      t2adda <= "11111010";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                  
                                  
                elsif cntr1 ="001100000100" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111011";
                      t2adda <= "11111011";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                        
                                        
                                        
                elsif cntr1 ="001100000101" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111100";
                      t2adda <= "11111100";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                                              
                                              
                elsif cntr1 ="001100000110" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111101";
                      t2adda <= "11111101";
                      t1dina <= bfrjout;
                      t2dina <= bfrjplout;
                                                    
                                                    
                                                    
                elsif cntr1 ="001100000111" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111110";
                      t2adda <= "11111110";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                                         
                                                         
                elsif cntr1 ="001100001000" THEN
                      
                      
                      t1wea <= '1';
                      t2wea <= '1';
                      t1adda <= "11111111";
                      t2adda <= "11111111";
                      t1dina <= bfrjplout;
                      t2dina <= bfrjout;
                                                             
                                                             
                                                             
                elsif cntr1 ="001100001001" THEN		
                
                
					  iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000000000";
                      ioaddb <= "000000010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100001010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000000001";
                      ioaddb <= "000000011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100001011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000000100";
                      ioaddb <= "000000110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100001100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000000101";
                      ioaddb <= "000000111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100001101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000001000";
                      ioaddb <= "000001010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100001110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000001001";
                      ioaddb <= "000001011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100001111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000001100";
                      ioaddb <= "000001110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100010000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000001101";
                      ioaddb <= "000001111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100010001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000010000";
                      ioaddb <= "000010010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100010010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000010001";
                      ioaddb <= "000010011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100010011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000010100";
                      ioaddb <= "000010110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100010100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000010101";
                      ioaddb <= "000010111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100010101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000011000";
                      ioaddb <= "000011010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100010110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000011001";
                      ioaddb <= "000011011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100010111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000011100";
                      ioaddb <= "000011110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100011000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000011101";
                      ioaddb <= "000011111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100011001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000100000";
                      ioaddb <= "000100010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100011010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000100001";
                      ioaddb <= "000100011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100011011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000100100";
                      ioaddb <= "000100110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100011100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000100101";
                      ioaddb <= "000100111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100011101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000101000";
                      ioaddb <= "000101010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100011110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000101001";
                      ioaddb <= "000101011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100011111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000101100";
                      ioaddb <= "000101110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100100000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000101101";
                      ioaddb <= "000101111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100100001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000110000";
                      ioaddb <= "000110010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100100010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000110001";
                      ioaddb <= "000110011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100100011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000110100";
                      ioaddb <= "000110110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100100100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000110101";
                      ioaddb <= "000110111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100100101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000111000";
                      ioaddb <= "000111010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100100110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000111001";
                      ioaddb <= "000111011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100100111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000111100";
                      ioaddb <= "000111110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100101000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "000111101";
                      ioaddb <= "000111111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100101001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001000000";
                      ioaddb <= "001000010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100101010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001000001";
                      ioaddb <= "001000011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100101011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001000100";
                      ioaddb <= "001000110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100101100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001000101";
                      ioaddb <= "001000111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100101101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001001000";
                      ioaddb <= "001001010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100101110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001001001";
                      ioaddb <= "001001011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100101111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001001100";
                      ioaddb <= "001001110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100110000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001001101";
                      ioaddb <= "001001111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100110001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001010000";
                      ioaddb <= "001010010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100110010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001010001";
                      ioaddb <= "001010011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100110011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001010100";
                      ioaddb <= "001010110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100110100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001010101";
                      ioaddb <= "001010111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100110101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001011000";
                      ioaddb <= "001011010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100110110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001011001";
                      ioaddb <= "001011011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100110111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001011100";
                      ioaddb <= "001011110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100111000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001011101";
                      ioaddb <= "001011111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100111001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001100000";
                      ioaddb <= "001100010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100111010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001100001";
                      ioaddb <= "001100011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100111011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001100100";
                      ioaddb <= "001100110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100111100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001100101";
                      ioaddb <= "001100111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100111101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001101000";
                      ioaddb <= "001101010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001100111110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001101001";
                      ioaddb <= "001101011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001100111111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001101100";
                      ioaddb <= "001101110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101000000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001101101";
                      ioaddb <= "001101111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101000001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001110000";
                      ioaddb <= "001110010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101000010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001110001";
                      ioaddb <= "001110011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101000011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001110100";
                      ioaddb <= "001110110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101000100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001110101";
                      ioaddb <= "001110111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101000101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001111000";
                      ioaddb <= "001111010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101000110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001111001";
                      ioaddb <= "001111011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101000111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001111100";
                      ioaddb <= "001111110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101001000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "001111101";
                      ioaddb <= "001111111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101001001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010000000";
                      ioaddb <= "010000010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101001010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010000001";
                      ioaddb <= "010000011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101001011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010000100";
                      ioaddb <= "010000110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101001100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010000101";
                      ioaddb <= "010000111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101001101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010001000";
                      ioaddb <= "010001010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101001110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010001001";
                      ioaddb <= "010001011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101001111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010001100";
                      ioaddb <= "010001110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101010000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010001101";
                      ioaddb <= "010001111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101010001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010010000";
                      ioaddb <= "010010010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101010010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010010001";
                      ioaddb <= "010010011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101010011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010010100";
                      ioaddb <= "010010110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101010100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010010101";
                      ioaddb <= "010010111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101010101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010011000";
                      ioaddb <= "010011010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101010110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010011001";
                      ioaddb <= "010011011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101010111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010011100";
                      ioaddb <= "010011110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101011000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010011101";
                      ioaddb <= "010011111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101011001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010100000";
                      ioaddb <= "010100010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101011010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010100001";
                      ioaddb <= "010100011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101011011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010100100";
                      ioaddb <= "010100110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101011100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010100101";
                      ioaddb <= "010100111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101011101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010101000";
                      ioaddb <= "010101010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101011110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010101001";
                      ioaddb <= "010101011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101011111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010101100";
                      ioaddb <= "010101110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101100000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010101101";
                      ioaddb <= "010101111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101100001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010110000";
                      ioaddb <= "010110010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101100010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010110001";
                      ioaddb <= "010110011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101100011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010110100";
                      ioaddb <= "010110110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101100100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010110101";
                      ioaddb <= "010110111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101100101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010111000";
                      ioaddb <= "010111010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101100110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010111001";
                      ioaddb <= "010111011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101100111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010111100";
                      ioaddb <= "010111110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101101000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "010111101";
                      ioaddb <= "010111111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101101001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011000000";
                      ioaddb <= "011000010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101101010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011000001";
                      ioaddb <= "011000011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101101011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011000100";
                      ioaddb <= "011000110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101101100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011000101";
                      ioaddb <= "011000111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101101101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011001000";
                      ioaddb <= "011001010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101101110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011001001";
                      ioaddb <= "011001011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101101111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011001100";
                      ioaddb <= "011001110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101110000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011001101";
                      ioaddb <= "011001111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101110001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011010000";
                      ioaddb <= "011010010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101110010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011010001";
                      ioaddb <= "011010011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101110011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011010100";
                      ioaddb <= "011010110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101110100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011010101";
                      ioaddb <= "011010111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101110101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011011000";
                      ioaddb <= "011011010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101110110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011011001";
                      ioaddb <= "011011011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101110111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011011100";
                      ioaddb <= "011011110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101111000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011011101";
                      ioaddb <= "011011111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101111001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011100000";
                      ioaddb <= "011100010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101111010" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011100001";
                      ioaddb <= "011100011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101111011" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011100100";
                      ioaddb <= "011100110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101111100" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011100101";
                      ioaddb <= "011100111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101111101" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011101000";
                      ioaddb <= "011101010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001101111110" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011101001";
                      ioaddb <= "011101011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                      
                elsif cntr1 ="001101111111" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011101100";
                      ioaddb <= "011101110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                elsif cntr1 ="001110000000" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011101101";
                      ioaddb <= "011101111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                       
				elsif cntr1 ="001110000001" THEN
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011110000";
                      ioaddb <= "011110010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                      
                      
                       
                elsif cntr1 ="001110000010" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011110001";
                      ioaddb <= "011110011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                            
                            
                             
                elsif cntr1 ="001110000011" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011110100";
                      ioaddb <= "011110110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                  
                                  
                                   
                elsif cntr1 ="001110000100" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011110101";
                      ioaddb <= "011110111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                        
                                        
                                         
                elsif cntr1 ="001110000101" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011111000";
                      ioaddb <= "011111010";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                               
                                               
                                                
                 elsif cntr1 ="001110000110" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011111001";
                      ioaddb <= "011111011";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                                     
                                                     
                                                      
                 elsif cntr1 ="001110000111" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011111100";
                      ioaddb <= "011111110";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                                           
                                                           
                                                           
                 elsif cntr1 ="001110001000" THEN
                      
                      
                      
                      
                      
                      iowea <= '1';
                      ioweb <= '1';
                      ioadda <= "011111101";
                      ioaddb <= "011111111";
                      iodina <= bfrjout;
                      iodinb <= bfrjplout;
                                                           
                       
					
                                                           									
                 elsif cntr1 ="001110001001" THEN
				
					
                 elsif cntr1 ="001110001010" THEN
				
				
				
				END IF;
				
				
				
				
			
			ELSIF cur_st = toinvntt THEN
				
				IF cntr ="000000000000" THEN
				      ioadda <= "000000000";
				      ioaddb <= "000000010";
				      
					  bfmod <= "10";
					  
					  
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000001";
				ELSIF cntr ="000000000001" THEN
				      ioadda <= "000000001";
				      ioaddb <= "000000011";
				      
					  
				
				
				
				
				
				
				
				
				
				
				
				       zetain   <="01111111";
				      cntr <= "000000000010";
				ELSIF cntr ="000000000010" THEN
				      ioadda <= "000000100";
				      ioaddb <= "000000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000011";
				ELSIF cntr ="000000000011" THEN
				      ioadda <= "000000101";
				      ioaddb <= "000000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				       zetain   <="01111110";
				      cntr <= "000000000100";
				ELSIF cntr ="000000000100" THEN
				      ioadda <= "000001000";
				      ioaddb <= "000001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000101";
				ELSIF cntr ="000000000101" THEN
				      ioadda <= "000001001";
				      ioaddb <= "000001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				       zetain   <="01111101";
				      cntr <= "000000000110";
				ELSIF cntr ="000000000110" THEN
				      ioadda <= "000001100";
				      ioaddb <= "000001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000111";
				ELSIF cntr ="000000000111" THEN
				      ioadda <= "000001101";
				      ioaddb <= "000001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				       zetain   <="01111100";
				      cntr <= "000000001000";
				ELSIF cntr ="000000001000" THEN
				      ioadda <= "000010000";
				      ioaddb <= "000010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
					  
				
				
				
				
				
				
				
				
				      cntr <= "000000001001";
				ELSIF cntr ="000000001001" THEN
				      ioadda <= "000010001";
				      ioaddb <= "000010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
					  
				
				
				      
				      
				       zetain   <="01111011";
				      cntr <= "000000001010";
				ELSIF cntr ="000000001010" THEN
				      ioadda <= "000010100";
				      ioaddb <= "000010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001011";
				ELSIF cntr ="000000001011" THEN
				      ioadda <= "000010101";
				      ioaddb <= "000010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01111010";
				      cntr <= "000000001100";
				ELSIF cntr ="000000001100" THEN
				      ioadda <= "000011000";
				      ioaddb <= "000011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001101";
				ELSIF cntr ="000000001101" THEN
				      ioadda <= "000011001";
				      ioaddb <= "000011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01111001";
				      cntr <= "000000001110";
				ELSIF cntr ="000000001110" THEN
				      ioadda <= "000011100";
				      ioaddb <= "000011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001111";
				ELSIF cntr ="000000001111" THEN
				      ioadda <= "000011101";
				      ioaddb <= "000011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01111000";
				      cntr <= "000000010000";
				ELSIF cntr ="000000010000" THEN
				      ioadda <= "000100000";
				      ioaddb <= "000100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010001";
				ELSIF cntr ="000000010001" THEN
				      ioadda <= "000100001";
				      ioaddb <= "000100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110111";
				      cntr <= "000000010010";
				ELSIF cntr ="000000010010" THEN
				      ioadda <= "000100100";
				      ioaddb <= "000100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010011";
				ELSIF cntr ="000000010011" THEN
				      ioadda <= "000100101";
				      ioaddb <= "000100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110110";
				      cntr <= "000000010100";
				ELSIF cntr ="000000010100" THEN
				      ioadda <= "000101000";
				      ioaddb <= "000101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010101";
				ELSIF cntr ="000000010101" THEN
				      ioadda <= "000101001";
				      ioaddb <= "000101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110101";
				      cntr <= "000000010110";
				ELSIF cntr ="000000010110" THEN
				      ioadda <= "000101100";
				      ioaddb <= "000101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010111";
				ELSIF cntr ="000000010111" THEN
				      ioadda <= "000101101";
				      ioaddb <= "000101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110100";
				      cntr <= "000000011000";
				ELSIF cntr ="000000011000" THEN
				      ioadda <= "000110000";
				      ioaddb <= "000110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011001";
				ELSIF cntr ="000000011001" THEN
				      ioadda <= "000110001";
				      ioaddb <= "000110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110011";
				      cntr <= "000000011010";
				ELSIF cntr ="000000011010" THEN
				      ioadda <= "000110100";
				      ioaddb <= "000110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011011";
				ELSIF cntr ="000000011011" THEN
				      ioadda <= "000110101";
				      ioaddb <= "000110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110010";
				      cntr <= "000000011100";
				ELSIF cntr ="000000011100" THEN
				      ioadda <= "000111000";
				      ioaddb <= "000111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011101";
				ELSIF cntr ="000000011101" THEN
				      ioadda <= "000111001";
				      ioaddb <= "000111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110001";
				      cntr <= "000000011110";
				ELSIF cntr ="000000011110" THEN
				      ioadda <= "000111100";
				      ioaddb <= "000111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011111";
				ELSIF cntr ="000000011111" THEN
				      ioadda <= "000111101";
				      ioaddb <= "000111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01110000";
				      cntr <= "000000100000";
				ELSIF cntr ="000000100000" THEN
				      ioadda <= "001000000";
				      ioaddb <= "001000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100001";
				ELSIF cntr ="000000100001" THEN
				      ioadda <= "001000001";
				      ioaddb <= "001000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101111";
				      cntr <= "000000100010";
				ELSIF cntr ="000000100010" THEN
				      ioadda <= "001000100";
				      ioaddb <= "001000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100011";
				ELSIF cntr ="000000100011" THEN
				      ioadda <= "001000101";
				      ioaddb <= "001000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101110";
				      cntr <= "000000100100";
				ELSIF cntr ="000000100100" THEN
				      ioadda <= "001001000";
				      ioaddb <= "001001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100101";
				ELSIF cntr ="000000100101" THEN
				      ioadda <= "001001001";
				      ioaddb <= "001001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101101";
				      cntr <= "000000100110";
				ELSIF cntr ="000000100110" THEN
				      ioadda <= "001001100";
				      ioaddb <= "001001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100111";
				ELSIF cntr ="000000100111" THEN
				      ioadda <= "001001101";
				      ioaddb <= "001001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101100";
				      cntr <= "000000101000";
				ELSIF cntr ="000000101000" THEN
				      ioadda <= "001010000";
				      ioaddb <= "001010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101001";
				ELSIF cntr ="000000101001" THEN
				      ioadda <= "001010001";
				      ioaddb <= "001010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101011";
				      cntr <= "000000101010";
				ELSIF cntr ="000000101010" THEN
				      ioadda <= "001010100";
				      ioaddb <= "001010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101011";
				ELSIF cntr ="000000101011" THEN
				      ioadda <= "001010101";
				      ioaddb <= "001010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101010";
				      cntr <= "000000101100";
				ELSIF cntr ="000000101100" THEN
				      ioadda <= "001011000";
				      ioaddb <= "001011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101101";
				ELSIF cntr ="000000101101" THEN
				      ioadda <= "001011001";
				      ioaddb <= "001011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101001";
				      cntr <= "000000101110";
				ELSIF cntr ="000000101110" THEN
				      ioadda <= "001011100";
				      ioaddb <= "001011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101111";
				ELSIF cntr ="000000101111" THEN
				      ioadda <= "001011101";
				      ioaddb <= "001011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01101000";
				      cntr <= "000000110000";
				ELSIF cntr ="000000110000" THEN
				      ioadda <= "001100000";
				      ioaddb <= "001100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110001";
				ELSIF cntr ="000000110001" THEN
				      ioadda <= "001100001";
				      ioaddb <= "001100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100111";
				      cntr <= "000000110010";
				ELSIF cntr ="000000110010" THEN
				      ioadda <= "001100100";
				      ioaddb <= "001100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110011";
				ELSIF cntr ="000000110011" THEN
				      ioadda <= "001100101";
				      ioaddb <= "001100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100110";
				      cntr <= "000000110100";
				ELSIF cntr ="000000110100" THEN
				      ioadda <= "001101000";
				      ioaddb <= "001101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110101";
				ELSIF cntr ="000000110101" THEN
				      ioadda <= "001101001";
				      ioaddb <= "001101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100101";
				      cntr <= "000000110110";
				ELSIF cntr ="000000110110" THEN
				      ioadda <= "001101100";
				      ioaddb <= "001101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110111";
				ELSIF cntr ="000000110111" THEN
				      ioadda <= "001101101";
				      ioaddb <= "001101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100100";
				      cntr <= "000000111000";
				ELSIF cntr ="000000111000" THEN
				      ioadda <= "001110000";
				      ioaddb <= "001110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111001";
				ELSIF cntr ="000000111001" THEN
				      ioadda <= "001110001";
				      ioaddb <= "001110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100011";
				      cntr <= "000000111010";
				ELSIF cntr ="000000111010" THEN
				      ioadda <= "001110100";
				      ioaddb <= "001110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111011";
				ELSIF cntr ="000000111011" THEN
				      ioadda <= "001110101";
				      ioaddb <= "001110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100010";
				      cntr <= "000000111100";
				ELSIF cntr ="000000111100" THEN
				      ioadda <= "001111000";
				      ioaddb <= "001111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111101";
				ELSIF cntr ="000000111101" THEN
				      ioadda <= "001111001";
				      ioaddb <= "001111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100001";
				      cntr <= "000000111110";
				ELSIF cntr ="000000111110" THEN
				      ioadda <= "001111100";
				      ioaddb <= "001111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111111";
				ELSIF cntr ="000000111111" THEN
				      ioadda <= "001111101";
				      ioaddb <= "001111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01100000";
				      cntr <= "000001000000";
				ELSIF cntr ="000001000000" THEN
				      ioadda <= "010000000";
				      ioaddb <= "010000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000001";
				ELSIF cntr ="000001000001" THEN
				      ioadda <= "010000001";
				      ioaddb <= "010000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011111";
				      cntr <= "000001000010";
				ELSIF cntr ="000001000010" THEN
				      ioadda <= "010000100";
				      ioaddb <= "010000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000011";
				ELSIF cntr ="000001000011" THEN
				      ioadda <= "010000101";
				      ioaddb <= "010000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011110";
				      cntr <= "000001000100";
				ELSIF cntr ="000001000100" THEN
				      ioadda <= "010001000";
				      ioaddb <= "010001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000101";
				ELSIF cntr ="000001000101" THEN
				      ioadda <= "010001001";
				      ioaddb <= "010001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011101";
				      cntr <= "000001000110";
				ELSIF cntr ="000001000110" THEN
				      ioadda <= "010001100";
				      ioaddb <= "010001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000111";
				ELSIF cntr ="000001000111" THEN
				      ioadda <= "010001101";
				      ioaddb <= "010001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011100";
				      cntr <= "000001001000";
				ELSIF cntr ="000001001000" THEN
				      ioadda <= "010010000";
				      ioaddb <= "010010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001001";
				ELSIF cntr ="000001001001" THEN
				      ioadda <= "010010001";
				      ioaddb <= "010010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011011";
				      cntr <= "000001001010";
				ELSIF cntr ="000001001010" THEN
				      ioadda <= "010010100";
				      ioaddb <= "010010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001011";
				ELSIF cntr ="000001001011" THEN
				      ioadda <= "010010101";
				      ioaddb <= "010010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011010";
				      cntr <= "000001001100";
				ELSIF cntr ="000001001100" THEN
				      ioadda <= "010011000";
				      ioaddb <= "010011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001101";
				ELSIF cntr ="000001001101" THEN
				      ioadda <= "010011001";
				      ioaddb <= "010011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011001";
				      cntr <= "000001001110";
				ELSIF cntr ="000001001110" THEN
				      ioadda <= "010011100";
				      ioaddb <= "010011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001111";
				ELSIF cntr ="000001001111" THEN
				      ioadda <= "010011101";
				      ioaddb <= "010011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01011000";
				      cntr <= "000001010000";
				ELSIF cntr ="000001010000" THEN
				      ioadda <= "010100000";
				      ioaddb <= "010100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010001";
				ELSIF cntr ="000001010001" THEN
				      ioadda <= "010100001";
				      ioaddb <= "010100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010111";
				      cntr <= "000001010010";
				ELSIF cntr ="000001010010" THEN
				      ioadda <= "010100100";
				      ioaddb <= "010100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010011";
				ELSIF cntr ="000001010011" THEN
				      ioadda <= "010100101";
				      ioaddb <= "010100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010110";
				      cntr <= "000001010100";
				ELSIF cntr ="000001010100" THEN
				      ioadda <= "010101000";
				      ioaddb <= "010101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010101";
				ELSIF cntr ="000001010101" THEN
				      ioadda <= "010101001";
				      ioaddb <= "010101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010101";
				      cntr <= "000001010110";
				ELSIF cntr ="000001010110" THEN
				      ioadda <= "010101100";
				      ioaddb <= "010101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010111";
				ELSIF cntr ="000001010111" THEN
				      ioadda <= "010101101";
				      ioaddb <= "010101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010100";
				      cntr <= "000001011000";
				ELSIF cntr ="000001011000" THEN
				      ioadda <= "010110000";
				      ioaddb <= "010110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011001";
				ELSIF cntr ="000001011001" THEN
				      ioadda <= "010110001";
				      ioaddb <= "010110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010011";
				      cntr <= "000001011010";
				ELSIF cntr ="000001011010" THEN
				      ioadda <= "010110100";
				      ioaddb <= "010110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011011";
				ELSIF cntr ="000001011011" THEN
				      ioadda <= "010110101";
				      ioaddb <= "010110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010010";
				      cntr <= "000001011100";
				ELSIF cntr ="000001011100" THEN
				      ioadda <= "010111000";
				      ioaddb <= "010111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011101";
				ELSIF cntr ="000001011101" THEN
				      ioadda <= "010111001";
				      ioaddb <= "010111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010001";
				      cntr <= "000001011110";
				ELSIF cntr ="000001011110" THEN
				      ioadda <= "010111100";
				      ioaddb <= "010111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011111";
				ELSIF cntr ="000001011111" THEN
				      ioadda <= "010111101";
				      ioaddb <= "010111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01010000";
				      cntr <= "000001100000";
				ELSIF cntr ="000001100000" THEN
				      ioadda <= "011000000";
				      ioaddb <= "011000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100001";
				ELSIF cntr ="000001100001" THEN
				      ioadda <= "011000001";
				      ioaddb <= "011000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001111";
				      cntr <= "000001100010";
				ELSIF cntr ="000001100010" THEN
				      ioadda <= "011000100";
				      ioaddb <= "011000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100011";
				ELSIF cntr ="000001100011" THEN
				      ioadda <= "011000101";
				      ioaddb <= "011000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001110";
				      cntr <= "000001100100";
				ELSIF cntr ="000001100100" THEN
				      ioadda <= "011001000";
				      ioaddb <= "011001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100101";
				ELSIF cntr ="000001100101" THEN
				      ioadda <= "011001001";
				      ioaddb <= "011001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001101";
				      cntr <= "000001100110";
				ELSIF cntr ="000001100110" THEN
				      ioadda <= "011001100";
				      ioaddb <= "011001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100111";
				ELSIF cntr ="000001100111" THEN
				      ioadda <= "011001101";
				      ioaddb <= "011001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001100";
				      cntr <= "000001101000";
				ELSIF cntr ="000001101000" THEN
				      ioadda <= "011010000";
				      ioaddb <= "011010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101001";
				ELSIF cntr ="000001101001" THEN
				      ioadda <= "011010001";
				      ioaddb <= "011010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001011";
				      cntr <= "000001101010";
				ELSIF cntr ="000001101010" THEN
				      ioadda <= "011010100";
				      ioaddb <= "011010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101011";
				ELSIF cntr ="000001101011" THEN
				      ioadda <= "011010101";
				      ioaddb <= "011010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001010";
				      cntr <= "000001101100";
				ELSIF cntr ="000001101100" THEN
				      ioadda <= "011011000";
				      ioaddb <= "011011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101101";
				ELSIF cntr ="000001101101" THEN
				      ioadda <= "011011001";
				      ioaddb <= "011011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001001";
				      cntr <= "000001101110";
				ELSIF cntr ="000001101110" THEN
				      ioadda <= "011011100";
				      ioaddb <= "011011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101111";
				ELSIF cntr ="000001101111" THEN
				      ioadda <= "011011101";
				      ioaddb <= "011011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01001000";
				      cntr <= "000001110000";
				ELSIF cntr ="000001110000" THEN
				      ioadda <= "011100000";
				      ioaddb <= "011100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110001";
				ELSIF cntr ="000001110001" THEN
				      ioadda <= "011100001";
				      ioaddb <= "011100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000111";
				      cntr <= "000001110010";
				ELSIF cntr ="000001110010" THEN
				      ioadda <= "011100100";
				      ioaddb <= "011100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110011";
				ELSIF cntr ="000001110011" THEN
				      ioadda <= "011100101";
				      ioaddb <= "011100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000110";
				      cntr <= "000001110100";
				ELSIF cntr ="000001110100" THEN
				      ioadda <= "011101000";
				      ioaddb <= "011101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110101";
				ELSIF cntr ="000001110101" THEN
				      ioadda <= "011101001";
				      ioaddb <= "011101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000101";
				      cntr <= "000001110110";
				ELSIF cntr ="000001110110" THEN
				      ioadda <= "011101100";
				      ioaddb <= "011101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110111";
				ELSIF cntr ="000001110111" THEN
				      ioadda <= "011101101";
				      ioaddb <= "011101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000100";
				      cntr <= "000001111000";
				ELSIF cntr ="000001111000" THEN
				      ioadda <= "011110000";
				      ioaddb <= "011110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111001";
				ELSIF cntr ="000001111001" THEN
				      ioadda <= "011110001";
				      ioaddb <= "011110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000011";
				      cntr <= "000001111010";
				ELSIF cntr ="000001111010" THEN
				      ioadda <= "011110100";
				      ioaddb <= "011110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111011";
				ELSIF cntr ="000001111011" THEN
				      ioadda <= "011110101";
				      ioaddb <= "011110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000010";
				      cntr <= "000001111100";
				ELSIF cntr ="000001111100" THEN
				      ioadda <= "011111000";
				      ioaddb <= "011111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111101";
				ELSIF cntr ="000001111101" THEN
				      ioadda <= "011111001";
				      ioaddb <= "011111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000001";
				      cntr <= "000001111110";
				ELSIF cntr ="000001111110" THEN
				      ioadda <= "011111100";
				      ioaddb <= "011111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111111";
				ELSIF cntr ="000001111111" THEN
				      ioadda <= "011111101";
				      ioaddb <= "011111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				       zetain   <="01000000";
				      cntr <= "000010000000";
				ELSIF cntr ="000010000000" THEN
				      t1addb <= "00000000";	  
				      t2addb <= "00000010";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010000001";
				ELSIF cntr ="000010000001" THEN
				      t1addb <= "00000001";	  
				      t2addb <= "00000011";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				        zetain   <="00111111";      
				      cntr <= "000010000010";
				ELSIF cntr ="000010000010" THEN
				      t1addb <= "00000010";      
				      t2addb <= "00000000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000010000011";      
				ELSIF cntr ="000010000011" THEN      
				      t1addb <= "00000011";      
				      t2addb <= "00000001";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000010000100";          
				ELSIF cntr ="000010000100" THEN        
				      t1addb <= "00000100";      
				      t2addb <= "00000110";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000010000101";          
				ELSIF cntr ="000010000101" THEN        
				      t1addb <= "00000101";      
				      t2addb <= "00000111";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                              
				                              
				        zetain   <="00111110";                              
				      cntr <= "000010000110";              
				ELSIF cntr ="000010000110" THEN            
				      t1addb <= "00000110";      
				      t2addb <= "00000100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000010000111";            
				ELSIF cntr ="000010000111" THEN          
				      t1addb <= "00000111";      
				      t2addb <= "00000101";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                          
				                                          
				                                          
				      cntr <= "000010001000";             
				ELSIF cntr ="000010001000" THEN           
				      t1addb <= "00001000";      
				      t2addb <= "00001010";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                                         
				                                         										
				                                   
				      cntr <= "000010001001";      
				ELSIF cntr ="000010001001" THEN    
				      t1addb <= "00001001";
				      t2addb <= "00001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				
				
				      
				      
				        zetain   <="00111101";
				      cntr <= "000010001010";
				elsif cntr ="000010001010" THEN
				      t1addb <= "00001010";
				      t2addb <= "00001000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001011";
				elsif cntr ="000010001011" THEN
				      t1addb <= "00001011";
				      t2addb <= "00001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001100";
				elsif cntr ="000010001100" THEN
				      t1addb <= "00001100";
				      t2addb <= "00001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001101";
				elsif cntr ="000010001101" THEN
				      t1addb <= "00001101";
				      t2addb <= "00001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00111100";
				      cntr <= "000010001110";
				elsif cntr ="000010001110" THEN
				      t1addb <= "00001110";
				      t2addb <= "00001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001111";
				elsif cntr ="000010001111" THEN
				      t1addb <= "00001111";
				      t2addb <= "00001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010000";
				elsif cntr ="000010010000" THEN
				      t1addb <= "00010000";
				      t2addb <= "00010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010001";
				elsif cntr ="000010010001" THEN
				      t1addb <= "00010001";
				      t2addb <= "00010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00111011";
				      cntr <= "000010010010";
				elsif cntr ="000010010010" THEN
				      t1addb <= "00010010";
				      t2addb <= "00010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010011";
				elsif cntr ="000010010011" THEN
				      t1addb <= "00010011";
				      t2addb <= "00010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010100";
				elsif cntr ="000010010100" THEN
				      t1addb <= "00010100";
				      t2addb <= "00010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010101";
				elsif cntr ="000010010101" THEN
				      t1addb <= "00010101";
				      t2addb <= "00010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00111010";
				      cntr <= "000010010110";
				elsif cntr ="000010010110" THEN
				      t1addb <= "00010110";
				      t2addb <= "00010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010111";
				elsif cntr ="000010010111" THEN
				      t1addb <= "00010111";
				      t2addb <= "00010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011000";
				elsif cntr ="000010011000" THEN
				      t1addb <= "00011000";
				      t2addb <= "00011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011001";
				elsif cntr ="000010011001" THEN
				      t1addb <= "00011001";
				      t2addb <= "00011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00111001";
				      cntr <= "000010011010";
				elsif cntr ="000010011010" THEN
				      t1addb <= "00011010";
				      t2addb <= "00011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011011";
				elsif cntr ="000010011011" THEN
				      t1addb <= "00011011";
				      t2addb <= "00011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011100";
				elsif cntr ="000010011100" THEN
				      t1addb <= "00011100";
				      t2addb <= "00011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011101";
				elsif cntr ="000010011101" THEN
				      t1addb <= "00011101";
				      t2addb <= "00011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00111000";
				      cntr <= "000010011110";
				elsif cntr ="000010011110" THEN
				      t1addb <= "00011110";
				      t2addb <= "00011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011111";
				elsif cntr ="000010011111" THEN
				      t1addb <= "00011111";
				      t2addb <= "00011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100000";
				elsif cntr ="000010100000" THEN
				      t1addb <= "00100000";
				      t2addb <= "00100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100001";
				elsif cntr ="000010100001" THEN
				      t1addb <= "00100001";
				      t2addb <= "00100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110111";
				      cntr <= "000010100010";
				elsif cntr ="000010100010" THEN
				      t1addb <= "00100010";
				      t2addb <= "00100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100011";
				elsif cntr ="000010100011" THEN
				      t1addb <= "00100011";
				      t2addb <= "00100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100100";
				elsif cntr ="000010100100" THEN
				      t1addb <= "00100100";
				      t2addb <= "00100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100101";
				elsif cntr ="000010100101" THEN
				      t1addb <= "00100101";
				      t2addb <= "00100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110110";
				      cntr <= "000010100110";
				elsif cntr ="000010100110" THEN
				      t1addb <= "00100110";
				      t2addb <= "00100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100111";
				elsif cntr ="000010100111" THEN
				      t1addb <= "00100111";
				      t2addb <= "00100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101000";
				elsif cntr ="000010101000" THEN
				      t1addb <= "00101000";
				      t2addb <= "00101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101001";
				elsif cntr ="000010101001" THEN
				      t1addb <= "00101001";
				      t2addb <= "00101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110101";
				      cntr <= "000010101010";
				elsif cntr ="000010101010" THEN
				      t1addb <= "00101010";
				      t2addb <= "00101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101011";
				elsif cntr ="000010101011" THEN
				      t1addb <= "00101011";
				      t2addb <= "00101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101100";
				elsif cntr ="000010101100" THEN
				      t1addb <= "00101100";
				      t2addb <= "00101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101101";
				elsif cntr ="000010101101" THEN
				      t1addb <= "00101101";
				      t2addb <= "00101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110100";
				      cntr <= "000010101110";
				elsif cntr ="000010101110" THEN
				      t1addb <= "00101110";
				      t2addb <= "00101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101111";
				elsif cntr ="000010101111" THEN
				      t1addb <= "00101111";
				      t2addb <= "00101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110000";
				elsif cntr ="000010110000" THEN
				      t1addb <= "00110000";
				      t2addb <= "00110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110001";
				elsif cntr ="000010110001" THEN
				      t1addb <= "00110001";
				      t2addb <= "00110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110011";
				      cntr <= "000010110010";
				elsif cntr ="000010110010" THEN
				      t1addb <= "00110010";
				      t2addb <= "00110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110011";
				elsif cntr ="000010110011" THEN
				      t1addb <= "00110011";
				      t2addb <= "00110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110100";
				elsif cntr ="000010110100" THEN
				      t1addb <= "00110100";
				      t2addb <= "00110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110101";
				elsif cntr ="000010110101" THEN
				      t1addb <= "00110101";
				      t2addb <= "00110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110010";
				      cntr <= "000010110110";
				elsif cntr ="000010110110" THEN
				      t1addb <= "00110110";
				      t2addb <= "00110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110111";
				elsif cntr ="000010110111" THEN
				      t1addb <= "00110111";
				      t2addb <= "00110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111000";
				elsif cntr ="000010111000" THEN
				      t1addb <= "00111000";
				      t2addb <= "00111010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111001";
				elsif cntr ="000010111001" THEN
				      t1addb <= "00111001";
				      t2addb <= "00111011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110001";
				      cntr <= "000010111010";
				elsif cntr ="000010111010" THEN
				      t1addb <= "00111010";
				      t2addb <= "00111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111011";
				elsif cntr ="000010111011" THEN
				      t1addb <= "00111011";
				      t2addb <= "00111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111100";
				elsif cntr ="000010111100" THEN
				      t1addb <= "00111100";
				      t2addb <= "00111110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111101";
				elsif cntr ="000010111101" THEN
				      t1addb <= "00111101";
				      t2addb <= "00111111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00110000";
				      cntr <= "000010111110";
				elsif cntr ="000010111110" THEN
				      t1addb <= "00111110";
				      t2addb <= "00111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111111";
				elsif cntr ="000010111111" THEN
				      t1addb <= "00111111";
				      t2addb <= "00111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000000";
				elsif cntr ="000011000000" THEN
				      t1addb <= "01000000";
				      t2addb <= "01000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000001";
				elsif cntr ="000011000001" THEN
				      t1addb <= "01000001";
				      t2addb <= "01000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101111";
				      cntr <= "000011000010";
				elsif cntr ="000011000010" THEN
				      t1addb <= "01000010";
				      t2addb <= "01000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000011";
				elsif cntr ="000011000011" THEN
				      t1addb <= "01000011";
				      t2addb <= "01000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000100";
				elsif cntr ="000011000100" THEN
				      t1addb <= "01000100";
				      t2addb <= "01000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000101";
				elsif cntr ="000011000101" THEN
				      t1addb <= "01000101";
				      t2addb <= "01000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101110";
				      cntr <= "000011000110";
				elsif cntr ="000011000110" THEN
				      t1addb <= "01000110";
				      t2addb <= "01000100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000111";
				elsif cntr ="000011000111" THEN
				      t1addb <= "01000111";
				      t2addb <= "01000101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001000";
				elsif cntr ="000011001000" THEN
				      t1addb <= "01001000";
				      t2addb <= "01001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001001";
				elsif cntr ="000011001001" THEN
				      t1addb <= "01001001";
				      t2addb <= "01001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101101";
				      cntr <= "000011001010";
				elsif cntr ="000011001010" THEN
				      t1addb <= "01001010";
				      t2addb <= "01001000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001011";
				elsif cntr ="000011001011" THEN
				      t1addb <= "01001011";
				      t2addb <= "01001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001100";
				elsif cntr ="000011001100" THEN
				      t1addb <= "01001100";
				      t2addb <= "01001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001101";
				elsif cntr ="000011001101" THEN
				      t1addb <= "01001101";
				      t2addb <= "01001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101100";
				      cntr <= "000011001110";
				elsif cntr ="000011001110" THEN
				      t1addb <= "01001110";
				      t2addb <= "01001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001111";
				elsif cntr ="000011001111" THEN
				      t1addb <= "01001111";
				      t2addb <= "01001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010000";
				elsif cntr ="000011010000" THEN
				      t1addb <= "01010000";
				      t2addb <= "01010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010001";
				elsif cntr ="000011010001" THEN
				      t1addb <= "01010001";
				      t2addb <= "01010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101011";
				      cntr <= "000011010010";
				elsif cntr ="000011010010" THEN
				      t1addb <= "01010010";
				      t2addb <= "01010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010011";
				elsif cntr ="000011010011" THEN
				      t1addb <= "01010011";
				      t2addb <= "01010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010100";
				elsif cntr ="000011010100" THEN
				      t1addb <= "01010100";
				      t2addb <= "01010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010101";
				elsif cntr ="000011010101" THEN
				      t1addb <= "01010101";
				      t2addb <= "01010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101010";
				      cntr <= "000011010110";
				elsif cntr ="000011010110" THEN
				      t1addb <= "01010110";
				      t2addb <= "01010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010111";
				elsif cntr ="000011010111" THEN
				      t1addb <= "01010111";
				      t2addb <= "01010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011000";
				elsif cntr ="000011011000" THEN
				      t1addb <= "01011000";
				      t2addb <= "01011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011001";
				elsif cntr ="000011011001" THEN
				      t1addb <= "01011001";
				      t2addb <= "01011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101001";
				      cntr <= "000011011010";
				elsif cntr ="000011011010" THEN
				      t1addb <= "01011010";
				      t2addb <= "01011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011011";
				elsif cntr ="000011011011" THEN
				      t1addb <= "01011011";
				      t2addb <= "01011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011100";
				elsif cntr ="000011011100" THEN
				      t1addb <= "01011100";
				      t2addb <= "01011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011101";
				elsif cntr ="000011011101" THEN
				      t1addb <= "01011101";
				      t2addb <= "01011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00101000";
				      cntr <= "000011011110";
				elsif cntr ="000011011110" THEN
				      t1addb <= "01011110";
				      t2addb <= "01011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011111";
				elsif cntr ="000011011111" THEN
				      t1addb <= "01011111";
				      t2addb <= "01011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100000";
				elsif cntr ="000011100000" THEN
				      t1addb <= "01100000";
				      t2addb <= "01100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100001";
				elsif cntr ="000011100001" THEN
				      t1addb <= "01100001";
				      t2addb <= "01100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100111";
				      cntr <= "000011100010";
				elsif cntr ="000011100010" THEN
				      t1addb <= "01100010";
				      t2addb <= "01100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100011";
				elsif cntr ="000011100011" THEN
				      t1addb <= "01100011";
				      t2addb <= "01100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100100";
				elsif cntr ="000011100100" THEN
				      t1addb <= "01100100";
				      t2addb <= "01100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100101";
				elsif cntr ="000011100101" THEN
				      t1addb <= "01100101";
				      t2addb <= "01100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100110";
				      cntr <= "000011100110";
				elsif cntr ="000011100110" THEN
				      t1addb <= "01100110";
				      t2addb <= "01100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100111";
				elsif cntr ="000011100111" THEN
				      t1addb <= "01100111";
				      t2addb <= "01100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101000";
				elsif cntr ="000011101000" THEN
				      t1addb <= "01101000";
				      t2addb <= "01101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101001";
				elsif cntr ="000011101001" THEN
				      t1addb <= "01101001";
				      t2addb <= "01101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100101";
				      cntr <= "000011101010";
				elsif cntr ="000011101010" THEN
				      t1addb <= "01101010";
				      t2addb <= "01101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101011";
				elsif cntr ="000011101011" THEN
				      t1addb <= "01101011";
				      t2addb <= "01101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101100";
				elsif cntr ="000011101100" THEN
				      t1addb <= "01101100";
				      t2addb <= "01101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101101";
				elsif cntr ="000011101101" THEN
				      t1addb <= "01101101";
				      t2addb <= "01101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100100";
				      cntr <= "000011101110";
				elsif cntr ="000011101110" THEN
				      t1addb <= "01101110";
				      t2addb <= "01101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101111";
				elsif cntr ="000011101111" THEN
				      t1addb <= "01101111";
				      t2addb <= "01101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110000";
				elsif cntr ="000011110000" THEN
				      t1addb <= "01110000";
				      t2addb <= "01110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110001";
				elsif cntr ="000011110001" THEN
				      t1addb <= "01110001";
				      t2addb <= "01110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100011";
				      cntr <= "000011110010";
				elsif cntr ="000011110010" THEN
				      t1addb <= "01110010";
				      t2addb <= "01110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110011";
				elsif cntr ="000011110011" THEN
				      t1addb <= "01110011";
				      t2addb <= "01110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110100";
				elsif cntr ="000011110100" THEN
				      t1addb <= "01110100";
				      t2addb <= "01110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110101";
				elsif cntr ="000011110101" THEN
				      t1addb <= "01110101";
				      t2addb <= "01110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100010";
				      cntr <= "000011110110";
				elsif cntr ="000011110110" THEN
				      t1addb <= "01110110";
				      t2addb <= "01110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110111";
				elsif cntr ="000011110111" THEN
				      t1addb <= "01110111";
				      t2addb <= "01110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111000";
				elsif cntr ="000011111000" THEN
				      t1addb <= "01111000";
				      t2addb <= "01111010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111001";
				elsif cntr ="000011111001" THEN
				      t1addb <= "01111001";
				      t2addb <= "01111011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100001";
				      cntr <= "000011111010";
				elsif cntr ="000011111010" THEN
				      t1addb <= "01111010";
				      t2addb <= "01111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111011";
				elsif cntr ="000011111011" THEN
				      t1addb <= "01111011";
				      t2addb <= "01111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111100";
				elsif cntr ="000011111100" THEN
				      t1addb <= "01111100";
				      t2addb <= "01111110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111101";
				elsif cntr ="000011111101" THEN
				      t1addb <= "01111101";
				      t2addb <= "01111111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00100000";
				      cntr <= "000011111110";
				elsif cntr ="000011111110" THEN
				      t1addb <= "01111110";
				      t2addb <= "01111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111111";
				elsif cntr ="000011111111" THEN
				      t1addb <= "01111111";
				      t2addb <= "01111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100000000";  
				elsif cntr ="000100000000" THEN												
				      t1addb <= "10000000";      
				      t2addb <= "10000100";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100000001";  
				elsif cntr ="000100000001" THEN		
				      t1addb <= "10000001";      
				      t2addb <= "10000101";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011111";      
				      cntr <= "000100000010";  
				elsif cntr ="000100000010" THEN		
				      t1addb <= "10000010";      
				      t2addb <= "10000110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000100000011";        
				elsif cntr ="000100000011" THEN		      
				      t1addb <= "10000011";      
				      t2addb <= "10000111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000100000100";             
				elsif cntr ="000100000100" THEN		      
				      t1addb <= "10000100";      
				      t2addb <= "10000000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000100000101";             
				elsif cntr ="000100000101" THEN		      
				      t1addb <= "10000101";      
				      t2addb <= "10000001";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "000100000110";             
				elsif cntr ="000100000110" THEN		      
				      t1addb <= "10000110";      
				      t2addb <= "10000010";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000100000111";             
				elsif cntr ="000100000111" THEN		      
				      t1addb <= "10000111";      
				      t2addb <= "10000011";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                                          
				                                          
				                                          
				      cntr <= "000100001000";              
				elsif cntr ="000100001000" THEN		       
				      t1addb <= "10001000";      
				      t2addb <= "10001100";      
				      bfrjin     <= t2doutb;      
				      bfrjplin <= t1doutb;      
				      
				      
				      
				                                
				                                
				                                
				      cntr <= "000100001001";   
				elsif cntr ="000100001001" THEN	
				      t1addb <= "10001001";
				      t2addb <= "10001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				
				
				
				      
				      
				        zetain   <="00011110";
				      cntr <= "000100001010";
				elsif cntr ="000100001010" THEN
				      t1addb <= "10001010";
				      t2addb <= "10001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001011";
				elsif cntr ="000100001011" THEN
				      t1addb <= "10001011";
				      t2addb <= "10001111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001100";
				elsif cntr ="000100001100" THEN
				      t1addb <= "10001100";
				      t2addb <= "10001000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001101";
				elsif cntr ="000100001101" THEN
				      t1addb <= "10001101";
				      t2addb <= "10001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001110";
				elsif cntr ="000100001110" THEN
				      t1addb <= "10001110";
				      t2addb <= "10001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001111";
				elsif cntr ="000100001111" THEN
				      t1addb <= "10001111";
				      t2addb <= "10001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010000";
				elsif cntr ="000100010000" THEN
				      t1addb <= "10010000";
				      t2addb <= "10010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010001";
				elsif cntr ="000100010001" THEN
				      t1addb <= "10010001";
				      t2addb <= "10010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011101";
				      cntr <= "000100010010";
				elsif cntr ="000100010010" THEN
				      t1addb <= "10010010";
				      t2addb <= "10010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010011";
				elsif cntr ="000100010011" THEN
				      t1addb <= "10010011";
				      t2addb <= "10010111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010100";
				elsif cntr ="000100010100" THEN
				      t1addb <= "10010100";
				      t2addb <= "10010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010101";
				elsif cntr ="000100010101" THEN
				      t1addb <= "10010101";
				      t2addb <= "10010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010110";
				elsif cntr ="000100010110" THEN
				      t1addb <= "10010110";
				      t2addb <= "10010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010111";
				elsif cntr ="000100010111" THEN
				      t1addb <= "10010111";
				      t2addb <= "10010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011000";
				elsif cntr ="000100011000" THEN
				      t1addb <= "10011000";
				      t2addb <= "10011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011001";
				elsif cntr ="000100011001" THEN
				      t1addb <= "10011001";
				      t2addb <= "10011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011100";
				      cntr <= "000100011010";
				elsif cntr ="000100011010" THEN
				      t1addb <= "10011010";
				      t2addb <= "10011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011011";
				elsif cntr ="000100011011" THEN
				      t1addb <= "10011011";
				      t2addb <= "10011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011100";
				elsif cntr ="000100011100" THEN
				      t1addb <= "10011100";
				      t2addb <= "10011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011101";
				elsif cntr ="000100011101" THEN
				      t1addb <= "10011101";
				      t2addb <= "10011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011110";
				elsif cntr ="000100011110" THEN
				      t1addb <= "10011110";
				      t2addb <= "10011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011111";
				elsif cntr ="000100011111" THEN
				      t1addb <= "10011111";
				      t2addb <= "10011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100000";
				elsif cntr ="000100100000" THEN
				      t1addb <= "10100000";
				      t2addb <= "10100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100001";
				elsif cntr ="000100100001" THEN
				      t1addb <= "10100001";
				      t2addb <= "10100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011011";
				      cntr <= "000100100010";
				elsif cntr ="000100100010" THEN
				      t1addb <= "10100010";
				      t2addb <= "10100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100011";
				elsif cntr ="000100100011" THEN
				      t1addb <= "10100011";
				      t2addb <= "10100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100100";
				elsif cntr ="000100100100" THEN
				      t1addb <= "10100100";
				      t2addb <= "10100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100101";
				elsif cntr ="000100100101" THEN
				      t1addb <= "10100101";
				      t2addb <= "10100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100110";
				elsif cntr ="000100100110" THEN
				      t1addb <= "10100110";
				      t2addb <= "10100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100111";
				elsif cntr ="000100100111" THEN
				      t1addb <= "10100111";
				      t2addb <= "10100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101000";
				elsif cntr ="000100101000" THEN
				      t1addb <= "10101000";
				      t2addb <= "10101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101001";
				elsif cntr ="000100101001" THEN
				      t1addb <= "10101001";
				      t2addb <= "10101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011010";
				      cntr <= "000100101010";
				elsif cntr ="000100101010" THEN
				      t1addb <= "10101010";
				      t2addb <= "10101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101011";
				elsif cntr ="000100101011" THEN
				      t1addb <= "10101011";
				      t2addb <= "10101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101100";
				elsif cntr ="000100101100" THEN
				      t1addb <= "10101100";
				      t2addb <= "10101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101101";
				elsif cntr ="000100101101" THEN
				      t1addb <= "10101101";
				      t2addb <= "10101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101110";
				elsif cntr ="000100101110" THEN
				      t1addb <= "10101110";
				      t2addb <= "10101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101111";
				elsif cntr ="000100101111" THEN
				      t1addb <= "10101111";
				      t2addb <= "10101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110000";
				elsif cntr ="000100110000" THEN
				      t1addb <= "10110000";
				      t2addb <= "10110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110001";
				elsif cntr ="000100110001" THEN
				      t1addb <= "10110001";
				      t2addb <= "10110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011001";
				      cntr <= "000100110010";
				elsif cntr ="000100110010" THEN
				      t1addb <= "10110010";
				      t2addb <= "10110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110011";
				elsif cntr ="000100110011" THEN
				      t1addb <= "10110011";
				      t2addb <= "10110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110100";
				elsif cntr ="000100110100" THEN
				      t1addb <= "10110100";
				      t2addb <= "10110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110101";
				elsif cntr ="000100110101" THEN
				      t1addb <= "10110101";
				      t2addb <= "10110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110110";
				elsif cntr ="000100110110" THEN
				      t1addb <= "10110110";
				      t2addb <= "10110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110111";
				elsif cntr ="000100110111" THEN
				      t1addb <= "10110111";
				      t2addb <= "10110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111000";
				elsif cntr ="000100111000" THEN
				      t1addb <= "10111000";
				      t2addb <= "10111100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111001";
				elsif cntr ="000100111001" THEN
				      t1addb <= "10111001";
				      t2addb <= "10111101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00011000";
				      cntr <= "000100111010";
				elsif cntr ="000100111010" THEN
				      t1addb <= "10111010";
				      t2addb <= "10111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111011";
				elsif cntr ="000100111011" THEN
				      t1addb <= "10111011";
				      t2addb <= "10111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111100";
				elsif cntr ="000100111100" THEN
				      t1addb <= "10111100";
				      t2addb <= "10111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111101";
				elsif cntr ="000100111101" THEN
				      t1addb <= "10111101";
				      t2addb <= "10111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111110";
				elsif cntr ="000100111110" THEN
				      t1addb <= "10111110";
				      t2addb <= "10111010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111111";
				elsif cntr ="000100111111" THEN
				      t1addb <= "10111111";
				      t2addb <= "10111011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000000";
				elsif cntr ="000101000000" THEN
				      t1addb <= "11000000";
				      t2addb <= "11000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000001";
				elsif cntr ="000101000001" THEN
				      t1addb <= "11000001";
				      t2addb <= "11000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010111";
				      cntr <= "000101000010";
				elsif cntr ="000101000010" THEN
				      t1addb <= "11000010";
				      t2addb <= "11000110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000011";
				elsif cntr ="000101000011" THEN
				      t1addb <= "11000011";
				      t2addb <= "11000111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000100";
				elsif cntr ="000101000100" THEN
				      t1addb <= "11000100";
				      t2addb <= "11000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000101";
				elsif cntr ="000101000101" THEN
				      t1addb <= "11000101";
				      t2addb <= "11000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000110";
				elsif cntr ="000101000110" THEN
				      t1addb <= "11000110";
				      t2addb <= "11000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000111";
				elsif cntr ="000101000111" THEN
				      t1addb <= "11000111";
				      t2addb <= "11000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001000";
				elsif cntr ="000101001000" THEN
				      t1addb <= "11001000";
				      t2addb <= "11001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001001";
				elsif cntr ="000101001001" THEN
				      t1addb <= "11001001";
				      t2addb <= "11001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010110";
				      cntr <= "000101001010";
				elsif cntr ="000101001010" THEN
				      t1addb <= "11001010";
				      t2addb <= "11001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001011";
				elsif cntr ="000101001011" THEN
				      t1addb <= "11001011";
				      t2addb <= "11001111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001100";
				elsif cntr ="000101001100" THEN
				      t1addb <= "11001100";
				      t2addb <= "11001000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001101";
				elsif cntr ="000101001101" THEN
				      t1addb <= "11001101";
				      t2addb <= "11001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001110";
				elsif cntr ="000101001110" THEN
				      t1addb <= "11001110";
				      t2addb <= "11001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001111";
				elsif cntr ="000101001111" THEN
				      t1addb <= "11001111";
				      t2addb <= "11001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010000";
				elsif cntr ="000101010000" THEN
				      t1addb <= "11010000";
				      t2addb <= "11010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010001";
				elsif cntr ="000101010001" THEN
				      t1addb <= "11010001";
				      t2addb <= "11010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010101";
				      cntr <= "000101010010";
				elsif cntr ="000101010010" THEN
				      t1addb <= "11010010";
				      t2addb <= "11010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010011";
				elsif cntr ="000101010011" THEN
				      t1addb <= "11010011";
				      t2addb <= "11010111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010100";
				elsif cntr ="000101010100" THEN
				      t1addb <= "11010100";
				      t2addb <= "11010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010101";
				elsif cntr ="000101010101" THEN
				      t1addb <= "11010101";
				      t2addb <= "11010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010110";
				elsif cntr ="000101010110" THEN
				      t1addb <= "11010110";
				      t2addb <= "11010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010111";
				elsif cntr ="000101010111" THEN
				      t1addb <= "11010111";
				      t2addb <= "11010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011000";
				elsif cntr ="000101011000" THEN
				      t1addb <= "11011000";
				      t2addb <= "11011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011001";
				elsif cntr ="000101011001" THEN
				      t1addb <= "11011001";
				      t2addb <= "11011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010100";
				      cntr <= "000101011010";
				elsif cntr ="000101011010" THEN
				      t1addb <= "11011010";
				      t2addb <= "11011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011011";
				elsif cntr ="000101011011" THEN
				      t1addb <= "11011011";
				      t2addb <= "11011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011100";
				elsif cntr ="000101011100" THEN
				      t1addb <= "11011100";
				      t2addb <= "11011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011101";
				elsif cntr ="000101011101" THEN
				      t1addb <= "11011101";
				      t2addb <= "11011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011110";
				elsif cntr ="000101011110" THEN
				      t1addb <= "11011110";
				      t2addb <= "11011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011111";
				elsif cntr ="000101011111" THEN
				      t1addb <= "11011111";
				      t2addb <= "11011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100000";
				elsif cntr ="000101100000" THEN
				      t1addb <= "11100000";
				      t2addb <= "11100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100001";
				elsif cntr ="000101100001" THEN
				      t1addb <= "11100001";
				      t2addb <= "11100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010011";
				      cntr <= "000101100010";
				elsif cntr ="000101100010" THEN
				      t1addb <= "11100010";
				      t2addb <= "11100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100011";
				elsif cntr ="000101100011" THEN
				      t1addb <= "11100011";
				      t2addb <= "11100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100100";
				elsif cntr ="000101100100" THEN
				      t1addb <= "11100100";
				      t2addb <= "11100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100101";
				elsif cntr ="000101100101" THEN
				      t1addb <= "11100101";
				      t2addb <= "11100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100110";
				elsif cntr ="000101100110" THEN
				      t1addb <= "11100110";
				      t2addb <= "11100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100111";
				elsif cntr ="000101100111" THEN
				      t1addb <= "11100111";
				      t2addb <= "11100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101000";
				elsif cntr ="000101101000" THEN
				      t1addb <= "11101000";
				      t2addb <= "11101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101001";
				elsif cntr ="000101101001" THEN
				      t1addb <= "11101001";
				      t2addb <= "11101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010010";
				      cntr <= "000101101010";
				elsif cntr ="000101101010" THEN
				      t1addb <= "11101010";
				      t2addb <= "11101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101011";
				elsif cntr ="000101101011" THEN
				      t1addb <= "11101011";
				      t2addb <= "11101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101100";
				elsif cntr ="000101101100" THEN
				      t1addb <= "11101100";
				      t2addb <= "11101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101101";
				elsif cntr ="000101101101" THEN
				      t1addb <= "11101101";
				      t2addb <= "11101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101110";
				elsif cntr ="000101101110" THEN
				      t1addb <= "11101110";
				      t2addb <= "11101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101111";
				elsif cntr ="000101101111" THEN
				      t1addb <= "11101111";
				      t2addb <= "11101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110000";
				elsif cntr ="000101110000" THEN
				      t1addb <= "11110000";
				      t2addb <= "11110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110001";
				elsif cntr ="000101110001" THEN
				      t1addb <= "11110001";
				      t2addb <= "11110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010001";
				      cntr <= "000101110010";
				elsif cntr ="000101110010" THEN
				      t1addb <= "11110010";
				      t2addb <= "11110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110011";
				elsif cntr ="000101110011" THEN
				      t1addb <= "11110011";
				      t2addb <= "11110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110100";
				elsif cntr ="000101110100" THEN
				      t1addb <= "11110100";
				      t2addb <= "11110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110101";
				elsif cntr ="000101110101" THEN
				      t1addb <= "11110101";
				      t2addb <= "11110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110110";
				elsif cntr ="000101110110" THEN
				      t1addb <= "11110110";
				      t2addb <= "11110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110111";
				elsif cntr ="000101110111" THEN
				      t1addb <= "11110111";
				      t2addb <= "11110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111000";
				elsif cntr ="000101111000" THEN
				      t1addb <= "11111000";
				      t2addb <= "11111100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111001";
				elsif cntr ="000101111001" THEN
				      t1addb <= "11111001";
				      t2addb <= "11111101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00010000";
				      cntr <= "000101111010";
				elsif cntr ="000101111010" THEN
				      t1addb <= "11111010";
				      t2addb <= "11111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111011";
				elsif cntr ="000101111011" THEN
				      t1addb <= "11111011";
				      t2addb <= "11111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111100";
				elsif cntr ="000101111100" THEN
				      t1addb <= "11111100";
				      t2addb <= "11111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111101";
				elsif cntr ="000101111101" THEN
				      t1addb <= "11111101";
				      t2addb <= "11111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111110";
				elsif cntr ="000101111110" THEN
				      t1addb <= "11111110";
				      t2addb <= "11111010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111111";
				elsif cntr ="000101111111" THEN
				      t1addb <= "11111111";
				      t2addb <= "11111011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110000000";
				elsif cntr ="000110000000" THEN											
				      t1addb <= "00000000";      
				      t2addb <= "00001000";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110000001";
				elsif cntr ="000110000001" THEN	
				      t1addb <= "00000001";      
				      t2addb <= "00001001";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001111";      
				      cntr <= "000110000010";
				elsif cntr ="000110000010" THEN	
				      t1addb <= "00000010";      
				      t2addb <= "00001010";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000110000011";      
				elsif cntr ="000110000011" THEN	      
				      t1addb <= "00000011";      
				      t2addb <= "00001011";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000110000100";            
				elsif cntr ="000110000100" THEN	            
				      t1addb <= "00000100";      
				      t2addb <= "00001100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000110000101";            
				elsif cntr ="000110000101" THEN	         
				      t1addb <= "00000101";      
				      t2addb <= "00001101";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "000110000110";           
				elsif cntr ="000110000110" THEN	        
				      t1addb <= "00000110";      
				      t2addb <= "00001110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000110000111";           
				elsif cntr ="000110000111" THEN	        
				      t1addb <= "00000111";      
				      t2addb <= "00001111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                        
				                                        
				                                        
				      cntr <= "000110001000";           
				elsif cntr ="000110001000" THEN	        
				      t1addb <= "00001000";      
				      t2addb <= "00000000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                      
				                                      
				                                      
				      cntr <= "000110001001";         
				elsif cntr ="000110001001" THEN	      									
				      t1addb <= "00001001";
				      t2addb <= "00000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "000110001010";
				elsif cntr ="000110001010" THEN
				      t1addb <= "00001010";
				      t2addb <= "00000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001011";
				elsif cntr ="000110001011" THEN
				      t1addb <= "00001011";
				      t2addb <= "00000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001100";
				elsif cntr ="000110001100" THEN
				      t1addb <= "00001100";
				      t2addb <= "00000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001101";
				elsif cntr ="000110001101" THEN
				      t1addb <= "00001101";
				      t2addb <= "00000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001110";
				elsif cntr ="000110001110" THEN
				      t1addb <= "00001110";
				      t2addb <= "00000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001111";
				elsif cntr ="000110001111" THEN
				      t1addb <= "00001111";
				      t2addb <= "00000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010000";
				elsif cntr ="000110010000" THEN
				      t1addb <= "00010000";
				      t2addb <= "00011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010001";
				elsif cntr ="000110010001" THEN
				      t1addb <= "00010001";
				      t2addb <= "00011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001110";
				      cntr <= "000110010010";
				elsif cntr ="000110010010" THEN
				      t1addb <= "00010010";
				      t2addb <= "00011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010011";
				elsif cntr ="000110010011" THEN
				      t1addb <= "00010011";
				      t2addb <= "00011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010100";
				elsif cntr ="000110010100" THEN
				      t1addb <= "00010100";
				      t2addb <= "00011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010101";
				elsif cntr ="000110010101" THEN
				      t1addb <= "00010101";
				      t2addb <= "00011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010110";
				elsif cntr ="000110010110" THEN
				      t1addb <= "00010110";
				      t2addb <= "00011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010111";
				elsif cntr ="000110010111" THEN
				      t1addb <= "00010111";
				      t2addb <= "00011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011000";
				elsif cntr ="000110011000" THEN
				      t1addb <= "00011000";
				      t2addb <= "00010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011001";
				elsif cntr ="000110011001" THEN
				      t1addb <= "00011001";
				      t2addb <= "00010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011010";
				elsif cntr ="000110011010" THEN
				      t1addb <= "00011010";
				      t2addb <= "00010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011011";
				elsif cntr ="000110011011" THEN
				      t1addb <= "00011011";
				      t2addb <= "00010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011100";
				elsif cntr ="000110011100" THEN
				      t1addb <= "00011100";
				      t2addb <= "00010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011101";
				elsif cntr ="000110011101" THEN
				      t1addb <= "00011101";
				      t2addb <= "00010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011110";
				elsif cntr ="000110011110" THEN
				      t1addb <= "00011110";
				      t2addb <= "00010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011111";
				elsif cntr ="000110011111" THEN
				      t1addb <= "00011111";
				      t2addb <= "00010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100000";
				elsif cntr ="000110100000" THEN
				      t1addb <= "00100000";
				      t2addb <= "00101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100001";
				elsif cntr ="000110100001" THEN
				      t1addb <= "00100001";
				      t2addb <= "00101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001101";
				      cntr <= "000110100010";
				elsif cntr ="000110100010" THEN
				      t1addb <= "00100010";
				      t2addb <= "00101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100011";
				elsif cntr ="000110100011" THEN
				      t1addb <= "00100011";
				      t2addb <= "00101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100100";
				elsif cntr ="000110100100" THEN
				      t1addb <= "00100100";
				      t2addb <= "00101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100101";
				elsif cntr ="000110100101" THEN
				      t1addb <= "00100101";
				      t2addb <= "00101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100110";
				elsif cntr ="000110100110" THEN
				      t1addb <= "00100110";
				      t2addb <= "00101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100111";
				elsif cntr ="000110100111" THEN
				      t1addb <= "00100111";
				      t2addb <= "00101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101000";
				elsif cntr ="000110101000" THEN
				      t1addb <= "00101000";
				      t2addb <= "00100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101001";
				elsif cntr ="000110101001" THEN
				      t1addb <= "00101001";
				      t2addb <= "00100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101010";
				elsif cntr ="000110101010" THEN
				      t1addb <= "00101010";
				      t2addb <= "00100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101011";
				elsif cntr ="000110101011" THEN
				      t1addb <= "00101011";
				      t2addb <= "00100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101100";
				elsif cntr ="000110101100" THEN
				      t1addb <= "00101100";
				      t2addb <= "00100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101101";
				elsif cntr ="000110101101" THEN
				      t1addb <= "00101101";
				      t2addb <= "00100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101110";
				elsif cntr ="000110101110" THEN
				      t1addb <= "00101110";
				      t2addb <= "00100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101111";
				elsif cntr ="000110101111" THEN
				      t1addb <= "00101111";
				      t2addb <= "00100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110000";
				elsif cntr ="000110110000" THEN
				      t1addb <= "00110000";
				      t2addb <= "00111000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110001";
				elsif cntr ="000110110001" THEN
				      t1addb <= "00110001";
				      t2addb <= "00111001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001100";
				      cntr <= "000110110010";
				elsif cntr ="000110110010" THEN
				      t1addb <= "00110010";
				      t2addb <= "00111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110011";
				elsif cntr ="000110110011" THEN
				      t1addb <= "00110011";
				      t2addb <= "00111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110100";
				elsif cntr ="000110110100" THEN
				      t1addb <= "00110100";
				      t2addb <= "00111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110101";
				elsif cntr ="000110110101" THEN
				      t1addb <= "00110101";
				      t2addb <= "00111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110110";
				elsif cntr ="000110110110" THEN
				      t1addb <= "00110110";
				      t2addb <= "00111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110111";
				elsif cntr ="000110110111" THEN
				      t1addb <= "00110111";
				      t2addb <= "00111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111000";
				elsif cntr ="000110111000" THEN
				      t1addb <= "00111000";
				      t2addb <= "00110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111001";
				elsif cntr ="000110111001" THEN
				      t1addb <= "00111001";
				      t2addb <= "00110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111010";
				elsif cntr ="000110111010" THEN
				      t1addb <= "00111010";
				      t2addb <= "00110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111011";
				elsif cntr ="000110111011" THEN
				      t1addb <= "00111011";
				      t2addb <= "00110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111100";
				elsif cntr ="000110111100" THEN
				      t1addb <= "00111100";
				      t2addb <= "00110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111101";
				elsif cntr ="000110111101" THEN
				      t1addb <= "00111101";
				      t2addb <= "00110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111110";
				elsif cntr ="000110111110" THEN
				      t1addb <= "00111110";
				      t2addb <= "00110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111111";
				elsif cntr ="000110111111" THEN
				      t1addb <= "00111111";
				      t2addb <= "00110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000000";
				elsif cntr ="000111000000" THEN
				      t1addb <= "01000000";
				      t2addb <= "01001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000001";
				elsif cntr ="000111000001" THEN
				      t1addb <= "01000001";
				      t2addb <= "01001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001011";
				      cntr <= "000111000010";
				elsif cntr ="000111000010" THEN
				      t1addb <= "01000010";
				      t2addb <= "01001010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000011";
				elsif cntr ="000111000011" THEN
				      t1addb <= "01000011";
				      t2addb <= "01001011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000100";
				elsif cntr ="000111000100" THEN
				      t1addb <= "01000100";
				      t2addb <= "01001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000101";
				elsif cntr ="000111000101" THEN
				      t1addb <= "01000101";
				      t2addb <= "01001101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000110";
				elsif cntr ="000111000110" THEN
				      t1addb <= "01000110";
				      t2addb <= "01001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000111";
				elsif cntr ="000111000111" THEN
				      t1addb <= "01000111";
				      t2addb <= "01001111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001000";
				elsif cntr ="000111001000" THEN
				      t1addb <= "01001000";
				      t2addb <= "01000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001001";
				elsif cntr ="000111001001" THEN
				      t1addb <= "01001001";
				      t2addb <= "01000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001010";
				elsif cntr ="000111001010" THEN
				      t1addb <= "01001010";
				      t2addb <= "01000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001011";
				elsif cntr ="000111001011" THEN
				      t1addb <= "01001011";
				      t2addb <= "01000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001100";
				elsif cntr ="000111001100" THEN
				      t1addb <= "01001100";
				      t2addb <= "01000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001101";
				elsif cntr ="000111001101" THEN
				      t1addb <= "01001101";
				      t2addb <= "01000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001110";
				elsif cntr ="000111001110" THEN
				      t1addb <= "01001110";
				      t2addb <= "01000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001111";
				elsif cntr ="000111001111" THEN
				      t1addb <= "01001111";
				      t2addb <= "01000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010000";
				elsif cntr ="000111010000" THEN
				      t1addb <= "01010000";
				      t2addb <= "01011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010001";
				elsif cntr ="000111010001" THEN
				      t1addb <= "01010001";
				      t2addb <= "01011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001010";
				      cntr <= "000111010010";
				elsif cntr ="000111010010" THEN
				      t1addb <= "01010010";
				      t2addb <= "01011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010011";
				elsif cntr ="000111010011" THEN
				      t1addb <= "01010011";
				      t2addb <= "01011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010100";
				elsif cntr ="000111010100" THEN
				      t1addb <= "01010100";
				      t2addb <= "01011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010101";
				elsif cntr ="000111010101" THEN
				      t1addb <= "01010101";
				      t2addb <= "01011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010110";
				elsif cntr ="000111010110" THEN
				      t1addb <= "01010110";
				      t2addb <= "01011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010111";
				elsif cntr ="000111010111" THEN
				      t1addb <= "01010111";
				      t2addb <= "01011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011000";
				elsif cntr ="000111011000" THEN
				      t1addb <= "01011000";
				      t2addb <= "01010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011001";
				elsif cntr ="000111011001" THEN
				      t1addb <= "01011001";
				      t2addb <= "01010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011010";
				elsif cntr ="000111011010" THEN
				      t1addb <= "01011010";
				      t2addb <= "01010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011011";
				elsif cntr ="000111011011" THEN
				      t1addb <= "01011011";
				      t2addb <= "01010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011100";
				elsif cntr ="000111011100" THEN
				      t1addb <= "01011100";
				      t2addb <= "01010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011101";
				elsif cntr ="000111011101" THEN
				      t1addb <= "01011101";
				      t2addb <= "01010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011110";
				elsif cntr ="000111011110" THEN
				      t1addb <= "01011110";
				      t2addb <= "01010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011111";
				elsif cntr ="000111011111" THEN
				      t1addb <= "01011111";
				      t2addb <= "01010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100000";
				elsif cntr ="000111100000" THEN
				      t1addb <= "01100000";
				      t2addb <= "01101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100001";
				elsif cntr ="000111100001" THEN
				      t1addb <= "01100001";
				      t2addb <= "01101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001001";
				      cntr <= "000111100010";
				elsif cntr ="000111100010" THEN
				      t1addb <= "01100010";
				      t2addb <= "01101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100011";
				elsif cntr ="000111100011" THEN
				      t1addb <= "01100011";
				      t2addb <= "01101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100100";
				elsif cntr ="000111100100" THEN
				      t1addb <= "01100100";
				      t2addb <= "01101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100101";
				elsif cntr ="000111100101" THEN
				      t1addb <= "01100101";
				      t2addb <= "01101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100110";
				elsif cntr ="000111100110" THEN
				      t1addb <= "01100110";
				      t2addb <= "01101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100111";
				elsif cntr ="000111100111" THEN
				      t1addb <= "01100111";
				      t2addb <= "01101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101000";
				elsif cntr ="000111101000" THEN
				      t1addb <= "01101000";
				      t2addb <= "01100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101001";
				elsif cntr ="000111101001" THEN
				      t1addb <= "01101001";
				      t2addb <= "01100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101010";
				elsif cntr ="000111101010" THEN
				      t1addb <= "01101010";
				      t2addb <= "01100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101011";
				elsif cntr ="000111101011" THEN
				      t1addb <= "01101011";
				      t2addb <= "01100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101100";
				elsif cntr ="000111101100" THEN
				      t1addb <= "01101100";
				      t2addb <= "01100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101101";
				elsif cntr ="000111101101" THEN
				      t1addb <= "01101101";
				      t2addb <= "01100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101110";
				elsif cntr ="000111101110" THEN
				      t1addb <= "01101110";
				      t2addb <= "01100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101111";
				elsif cntr ="000111101111" THEN
				      t1addb <= "01101111";
				      t2addb <= "01100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110000";
				elsif cntr ="000111110000" THEN
				      t1addb <= "01110000";
				      t2addb <= "01111000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110001";
				elsif cntr ="000111110001" THEN
				      t1addb <= "01110001";
				      t2addb <= "01111001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00001000";
				      cntr <= "000111110010";
				elsif cntr ="000111110010" THEN
				      t1addb <= "01110010";
				      t2addb <= "01111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110011";
				elsif cntr ="000111110011" THEN
				      t1addb <= "01110011";
				      t2addb <= "01111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110100";
				elsif cntr ="000111110100" THEN
				      t1addb <= "01110100";
				      t2addb <= "01111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110101";
				elsif cntr ="000111110101" THEN
				      t1addb <= "01110101";
				      t2addb <= "01111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110110";
				elsif cntr ="000111110110" THEN
				      t1addb <= "01110110";
				      t2addb <= "01111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110111";
				elsif cntr ="000111110111" THEN
				      t1addb <= "01110111";
				      t2addb <= "01111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111000";
				elsif cntr ="000111111000" THEN
				      t1addb <= "01111000";
				      t2addb <= "01110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111001";
				elsif cntr ="000111111001" THEN
				      t1addb <= "01111001";
				      t2addb <= "01110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111010";
				elsif cntr ="000111111010" THEN
				      t1addb <= "01111010";
				      t2addb <= "01110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111011";
				elsif cntr ="000111111011" THEN
				      t1addb <= "01111011";
				      t2addb <= "01110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111100";
				elsif cntr ="000111111100" THEN
				      t1addb <= "01111100";
				      t2addb <= "01110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111101";
				elsif cntr ="000111111101" THEN
				      t1addb <= "01111101";
				      t2addb <= "01110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111110";
				elsif cntr ="000111111110" THEN
				      t1addb <= "01111110";
				      t2addb <= "01110110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111111";
				elsif cntr ="000111111111" THEN
				      t1addb <= "01111111";
				      t2addb <= "01110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000000000";				
				elsif cntr ="001000000000" THEN
				      t1addb <= "10000000";      
				      t2addb <= "10010000";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000000001";	
				elsif cntr ="001000000001" THEN
				      t1addb <= "10000001";      
				      t2addb <= "10010001";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000111";      
				      cntr <= "001000000010";	
				elsif cntr ="001000000010" THEN
				      t1addb <= "10000010";      
				      t2addb <= "10010010";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "001000000011";	      
				elsif cntr ="001000000011" THEN      
				      t1addb <= "10000011";      
				      t2addb <= "10010011";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001000000100";	       
				elsif cntr ="001000000100" THEN        
				      t1addb <= "10000100";      
				      t2addb <= "10010100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001000000101";	         
				elsif cntr ="001000000101" THEN          
				      t1addb <= "10000101";      
				      t2addb <= "10010101";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001000000110";	        
				elsif cntr ="001000000110" THEN         
				      t1addb <= "10000110";      
				      t2addb <= "10010110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001000000111";	          
				elsif cntr ="001000000111" THEN           
				      t1addb <= "10000111";      
				      t2addb <= "10010111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                         
				                                         
				                                         
				      cntr <= "001000001000";	         
				elsif cntr ="001000001000" THEN          
				      t1addb <= "10001000";      
				      t2addb <= "10011000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                  
				                                  
				                                  
				      cntr <= "001000001001";	  
				elsif cntr ="001000001001" THEN   
				      t1addb <= "10001001";
				      t2addb <= "10011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "001000001010";
				elsif cntr ="001000001010" THEN
				      t1addb <= "10001010";
				      t2addb <= "10011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001011";
				elsif cntr ="001000001011" THEN
				      t1addb <= "10001011";
				      t2addb <= "10011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001100";
				elsif cntr ="001000001100" THEN
				      t1addb <= "10001100";
				      t2addb <= "10011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001101";
				elsif cntr ="001000001101" THEN
				      t1addb <= "10001101";
				      t2addb <= "10011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001110";
				elsif cntr ="001000001110" THEN
				      t1addb <= "10001110";
				      t2addb <= "10011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001111";
				elsif cntr ="001000001111" THEN
				      t1addb <= "10001111";
				      t2addb <= "10011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010000";
				elsif cntr ="001000010000" THEN
				      t1addb <= "10010000";
				      t2addb <= "10000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010001";
				elsif cntr ="001000010001" THEN
				      t1addb <= "10010001";
				      t2addb <= "10000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010010";
				elsif cntr ="001000010010" THEN
				      t1addb <= "10010010";
				      t2addb <= "10000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010011";
				elsif cntr ="001000010011" THEN
				      t1addb <= "10010011";
				      t2addb <= "10000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010100";
				elsif cntr ="001000010100" THEN
				      t1addb <= "10010100";
				      t2addb <= "10000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010101";
				elsif cntr ="001000010101" THEN
				      t1addb <= "10010101";
				      t2addb <= "10000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010110";
				elsif cntr ="001000010110" THEN
				      t1addb <= "10010110";
				      t2addb <= "10000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010111";
				elsif cntr ="001000010111" THEN
				      t1addb <= "10010111";
				      t2addb <= "10000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011000";
				elsif cntr ="001000011000" THEN
				      t1addb <= "10011000";
				      t2addb <= "10001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011001";
				elsif cntr ="001000011001" THEN
				      t1addb <= "10011001";
				      t2addb <= "10001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011010";
				elsif cntr ="001000011010" THEN
				      t1addb <= "10011010";
				      t2addb <= "10001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011011";
				elsif cntr ="001000011011" THEN
				      t1addb <= "10011011";
				      t2addb <= "10001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011100";
				elsif cntr ="001000011100" THEN
				      t1addb <= "10011100";
				      t2addb <= "10001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011101";
				elsif cntr ="001000011101" THEN
				      t1addb <= "10011101";
				      t2addb <= "10001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011110";
				elsif cntr ="001000011110" THEN
				      t1addb <= "10011110";
				      t2addb <= "10001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011111";
				elsif cntr ="001000011111" THEN
				      t1addb <= "10011111";
				      t2addb <= "10001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100000";
				elsif cntr ="001000100000" THEN
				      t1addb <= "10100000";
				      t2addb <= "10110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100001";
				elsif cntr ="001000100001" THEN
				      t1addb <= "10100001";
				      t2addb <= "10110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000110";
				      cntr <= "001000100010";
				elsif cntr ="001000100010" THEN
				      t1addb <= "10100010";
				      t2addb <= "10110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100011";
				elsif cntr ="001000100011" THEN
				      t1addb <= "10100011";
				      t2addb <= "10110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100100";
				elsif cntr ="001000100100" THEN
				      t1addb <= "10100100";
				      t2addb <= "10110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100101";
				elsif cntr ="001000100101" THEN
				      t1addb <= "10100101";
				      t2addb <= "10110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100110";
				elsif cntr ="001000100110" THEN
				      t1addb <= "10100110";
				      t2addb <= "10110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100111";
				elsif cntr ="001000100111" THEN
				      t1addb <= "10100111";
				      t2addb <= "10110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101000";
				elsif cntr ="001000101000" THEN
				      t1addb <= "10101000";
				      t2addb <= "10111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101001";
				elsif cntr ="001000101001" THEN
				      t1addb <= "10101001";
				      t2addb <= "10111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101010";
				elsif cntr ="001000101010" THEN
				      t1addb <= "10101010";
				      t2addb <= "10111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101011";
				elsif cntr ="001000101011" THEN
				      t1addb <= "10101011";
				      t2addb <= "10111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101100";
				elsif cntr ="001000101100" THEN
				      t1addb <= "10101100";
				      t2addb <= "10111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101101";
				elsif cntr ="001000101101" THEN
				      t1addb <= "10101101";
				      t2addb <= "10111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101110";
				elsif cntr ="001000101110" THEN
				      t1addb <= "10101110";
				      t2addb <= "10111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101111";
				elsif cntr ="001000101111" THEN
				      t1addb <= "10101111";
				      t2addb <= "10111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110000";
				elsif cntr ="001000110000" THEN
				      t1addb <= "10110000";
				      t2addb <= "10100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110001";
				elsif cntr ="001000110001" THEN
				      t1addb <= "10110001";
				      t2addb <= "10100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110010";
				elsif cntr ="001000110010" THEN
				      t1addb <= "10110010";
				      t2addb <= "10100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110011";
				elsif cntr ="001000110011" THEN
				      t1addb <= "10110011";
				      t2addb <= "10100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110100";
				elsif cntr ="001000110100" THEN
				      t1addb <= "10110100";
				      t2addb <= "10100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110101";
				elsif cntr ="001000110101" THEN
				      t1addb <= "10110101";
				      t2addb <= "10100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110110";
				elsif cntr ="001000110110" THEN
				      t1addb <= "10110110";
				      t2addb <= "10100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110111";
				elsif cntr ="001000110111" THEN
				      t1addb <= "10110111";
				      t2addb <= "10100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111000";
				elsif cntr ="001000111000" THEN
				      t1addb <= "10111000";
				      t2addb <= "10101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111001";
				elsif cntr ="001000111001" THEN
				      t1addb <= "10111001";
				      t2addb <= "10101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111010";
				elsif cntr ="001000111010" THEN
				      t1addb <= "10111010";
				      t2addb <= "10101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111011";
				elsif cntr ="001000111011" THEN
				      t1addb <= "10111011";
				      t2addb <= "10101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111100";
				elsif cntr ="001000111100" THEN
				      t1addb <= "10111100";
				      t2addb <= "10101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111101";
				elsif cntr ="001000111101" THEN
				      t1addb <= "10111101";
				      t2addb <= "10101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111110";
				elsif cntr ="001000111110" THEN
				      t1addb <= "10111110";
				      t2addb <= "10101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111111";
				elsif cntr ="001000111111" THEN
				      t1addb <= "10111111";
				      t2addb <= "10101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000000";
				elsif cntr ="001001000000" THEN
				      t1addb <= "11000000";
				      t2addb <= "11010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000001";
				elsif cntr ="001001000001" THEN
				      t1addb <= "11000001";
				      t2addb <= "11010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000101";
				      cntr <= "001001000010";
				elsif cntr ="001001000010" THEN
				      t1addb <= "11000010";
				      t2addb <= "11010010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000011";
				elsif cntr ="001001000011" THEN
				      t1addb <= "11000011";
				      t2addb <= "11010011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000100";
				elsif cntr ="001001000100" THEN
				      t1addb <= "11000100";
				      t2addb <= "11010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000101";
				elsif cntr ="001001000101" THEN
				      t1addb <= "11000101";
				      t2addb <= "11010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000110";
				elsif cntr ="001001000110" THEN
				      t1addb <= "11000110";
				      t2addb <= "11010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000111";
				elsif cntr ="001001000111" THEN
				      t1addb <= "11000111";
				      t2addb <= "11010111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001000";
				elsif cntr ="001001001000" THEN
				      t1addb <= "11001000";
				      t2addb <= "11011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001001";
				elsif cntr ="001001001001" THEN
				      t1addb <= "11001001";
				      t2addb <= "11011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001010";
				elsif cntr ="001001001010" THEN
				      t1addb <= "11001010";
				      t2addb <= "11011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001011";
				elsif cntr ="001001001011" THEN
				      t1addb <= "11001011";
				      t2addb <= "11011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001100";
				elsif cntr ="001001001100" THEN
				      t1addb <= "11001100";
				      t2addb <= "11011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001101";
				elsif cntr ="001001001101" THEN
				      t1addb <= "11001101";
				      t2addb <= "11011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001110";
				elsif cntr ="001001001110" THEN
				      t1addb <= "11001110";
				      t2addb <= "11011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001111";
				elsif cntr ="001001001111" THEN
				      t1addb <= "11001111";
				      t2addb <= "11011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010000";
				elsif cntr ="001001010000" THEN
				      t1addb <= "11010000";
				      t2addb <= "11000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010001";
				elsif cntr ="001001010001" THEN
				      t1addb <= "11010001";
				      t2addb <= "11000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010010";
				elsif cntr ="001001010010" THEN
				      t1addb <= "11010010";
				      t2addb <= "11000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010011";
				elsif cntr ="001001010011" THEN
				      t1addb <= "11010011";
				      t2addb <= "11000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010100";
				elsif cntr ="001001010100" THEN
				      t1addb <= "11010100";
				      t2addb <= "11000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010101";
				elsif cntr ="001001010101" THEN
				      t1addb <= "11010101";
				      t2addb <= "11000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010110";
				elsif cntr ="001001010110" THEN
				      t1addb <= "11010110";
				      t2addb <= "11000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010111";
				elsif cntr ="001001010111" THEN
				      t1addb <= "11010111";
				      t2addb <= "11000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011000";
				elsif cntr ="001001011000" THEN
				      t1addb <= "11011000";
				      t2addb <= "11001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011001";
				elsif cntr ="001001011001" THEN
				      t1addb <= "11011001";
				      t2addb <= "11001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011010";
				elsif cntr ="001001011010" THEN
				      t1addb <= "11011010";
				      t2addb <= "11001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011011";
				elsif cntr ="001001011011" THEN
				      t1addb <= "11011011";
				      t2addb <= "11001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011100";
				elsif cntr ="001001011100" THEN
				      t1addb <= "11011100";
				      t2addb <= "11001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011101";
				elsif cntr ="001001011101" THEN
				      t1addb <= "11011101";
				      t2addb <= "11001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011110";
				elsif cntr ="001001011110" THEN
				      t1addb <= "11011110";
				      t2addb <= "11001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011111";
				elsif cntr ="001001011111" THEN
				      t1addb <= "11011111";
				      t2addb <= "11001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100000";
				elsif cntr ="001001100000" THEN
				      t1addb <= "11100000";
				      t2addb <= "11110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
						
				      
				      
				      
				      
				      
				      cntr <= "001001100001";
				elsif cntr ="001001100001" THEN
				      t1addb <= "11100001";
				      t2addb <= "11110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000100";
				      cntr <= "001001100010";
				elsif cntr ="001001100010" THEN
				      t1addb <= "11100010";
				      t2addb <= "11110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100011";
				elsif cntr ="001001100011" THEN
				      t1addb <= "11100011";
				      t2addb <= "11110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100100";
				elsif cntr ="001001100100" THEN
				      t1addb <= "11100100";
				      t2addb <= "11110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100101";
				elsif cntr ="001001100101" THEN
				      t1addb <= "11100101";
				      t2addb <= "11110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100110";
				elsif cntr ="001001100110" THEN
				      t1addb <= "11100110";
				      t2addb <= "11110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100111";
				elsif cntr ="001001100111" THEN
				      t1addb <= "11100111";		
				      t2addb <= "11110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101000";
				elsif cntr ="001001101000" THEN
				      t1addb <= "11101000";
				      t2addb <= "11111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101001";
				elsif cntr ="001001101001" THEN
				      t1addb <= "11101001";
				      t2addb <= "11111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101010";
				elsif cntr ="001001101010" THEN
				      t1addb <= "11101010";
				      t2addb <= "11111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101011";
				elsif cntr ="001001101011" THEN
				      t1addb <= "11101011";
				      t2addb <= "11111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101100";
				elsif cntr ="001001101100" THEN
				      t1addb <= "11101100";
				      t2addb <= "11111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101101";
				elsif cntr ="001001101101" THEN
				      t1addb <= "11101101";
				      t2addb <= "11111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
						
				      
				      cntr <= "001001101110";
				elsif cntr ="001001101110" THEN
				      t1addb <= "11101110";
				      t2addb <= "11111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101111";
				elsif cntr ="001001101111" THEN
				      t1addb <= "11101111";
				      t2addb <= "11111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110000";
				elsif cntr ="001001110000" THEN
				      t1addb <= "11110000";
				      t2addb <= "11100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110001";
				elsif cntr ="001001110001" THEN
				      t1addb <= "11110001";
				      t2addb <= "11100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;		
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110010";
				elsif cntr ="001001110010" THEN
				      t1addb <= "11110010";
				      t2addb <= "11100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110011";
				elsif cntr ="001001110011" THEN
				      t1addb <= "11110011";
				      t2addb <= "11100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110100";
				elsif cntr ="001001110100" THEN
				      t1addb <= "11110100";
				      t2addb <= "11100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110101";
				elsif cntr ="001001110101" THEN
				      t1addb <= "11110101";
				      t2addb <= "11100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110110";
				elsif cntr ="001001110110" THEN
				      t1addb <= "11110110";
				      t2addb <= "11100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110111";
				elsif cntr ="001001110111" THEN
				      t1addb <= "11110111";
				      t2addb <= "11100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111000";
				elsif cntr ="001001111000" THEN		
				      t1addb <= "11111000";
				      t2addb <= "11101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111001";
				elsif cntr ="001001111001" THEN
				      t1addb <= "11111001";
				      t2addb <= "11101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111010";
				elsif cntr ="001001111010" THEN
				      t1addb <= "11111010";
				      t2addb <= "11101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111011";
				elsif cntr ="001001111011" THEN
				      t1addb <= "11111011";
				      t2addb <= "11101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
						
				      
				      
				      
				      cntr <= "001001111100";
				elsif cntr ="001001111100" THEN
				      t1addb <= "11111100";
				      t2addb <= "11101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111101";
				elsif cntr ="001001111101" THEN
				      t1addb <= "11111101";
				      t2addb <= "11101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111110";
				elsif cntr ="001001111110" THEN
				      t1addb <= "11111110";
				      t2addb <= "11101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
						
				      
				      
				      cntr <= "001001111111";
				elsif cntr ="001001111111" THEN
				      t1addb <= "11111111";
				      t2addb <= "11101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010000000";
				elsif cntr ="001010000000" THEN												
				      t1addb <= "00000000";      
				      t2addb <= "00100000";      
				         bfrjin     <= t2doutb;
				         bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010000001";
				elsif cntr ="001010000001" THEN	
				      t1addb <= "00000001";      
				      t2addb <= "00100001";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000011";      
				      cntr <= "001010000010";
				elsif cntr ="001010000010" THEN	
				      t1addb <= "00000010";      
				      t2addb <= "00100010";      
				      bfrjin     <= t1doutb;		
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "001010000011";      
				elsif cntr ="001010000011" THEN	      
				      t1addb <= "00000011";      
				      t2addb <= "00100011";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001010000100";           
				elsif cntr ="001010000100" THEN	        
				      t1addb <= "00000100";      
				      t2addb <= "00100100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001010000101";           
				elsif cntr ="001010000101" THEN	        
				      t1addb <= "00000101";      
				      t2addb <= "00100101";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001010000110";         
				elsif cntr ="001010000110" THEN	      
				      t1addb <= "00000110";      
				      t2addb <= "00100110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001010000111";            
				elsif cntr ="001010000111" THEN	         
				      t1addb <= "00000111";      
				      t2addb <= "00100111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                       
				                                       
				                                       
				      cntr <= "001010001000";          
				elsif cntr ="001010001000" THEN	       
				      t1addb <= "00001000";      
				      t2addb <= "00101000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                         
				                                         
				                                         
				      cntr <= "001010001001";      											
				elsif cntr ="001010001001" THEN	   
				      t1addb <= "00001001";
				      t2addb <= "00101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "001010001010";
				elsif cntr ="001010001010" THEN
				      t1addb <= "00001010";
				      t2addb <= "00101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001011";
				elsif cntr ="001010001011" THEN
				      t1addb <= "00001011";
				      t2addb <= "00101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001100";
				elsif cntr ="001010001100" THEN
				      t1addb <= "00001100";
				      t2addb <= "00101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
						
				      
				      
				      
				      
				      cntr <= "001010001101";
				elsif cntr ="001010001101" THEN
				      t1addb <= "00001101";
				      t2addb <= "00101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001110";
				elsif cntr ="001010001110" THEN
				      t1addb <= "00001110";
				      t2addb <= "00101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001111";
				elsif cntr ="001010001111" THEN
				      t1addb <= "00001111";
				      t2addb <= "00101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010000";
				elsif cntr ="001010010000" THEN
				      t1addb <= "00010000";
				      t2addb <= "00110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010001";
				elsif cntr ="001010010001" THEN
				      t1addb <= "00010001";
				      t2addb <= "00110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010010";
				elsif cntr ="001010010010" THEN
				      t1addb <= "00010010";
				      t2addb <= "00110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010011";
				elsif cntr ="001010010011" THEN
				      t1addb <= "00010011";
				      t2addb <= "00110011";		
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010100";
				elsif cntr ="001010010100" THEN
				      t1addb <= "00010100";
				      t2addb <= "00110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010101";
				elsif cntr ="001010010101" THEN
				      t1addb <= "00010101";
				      t2addb <= "00110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010110";
				elsif cntr ="001010010110" THEN
				      t1addb <= "00010110";
				      t2addb <= "00110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010111";
				elsif cntr ="001010010111" THEN
				      t1addb <= "00010111";
				      t2addb <= "00110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011000";
				elsif cntr ="001010011000" THEN
				      t1addb <= "00011000";
				      t2addb <= "00111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011001";
				elsif cntr ="001010011001" THEN
				      t1addb <= "00011001";
				      t2addb <= "00111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
						
				      cntr <= "001010011010";
				elsif cntr ="001010011010" THEN
				      t1addb <= "00011010";
				      t2addb <= "00111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011011";
				elsif cntr ="001010011011" THEN
				      t1addb <= "00011011";
				      t2addb <= "00111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011100";
				elsif cntr ="001010011100" THEN
				      t1addb <= "00011100";
				      t2addb <= "00111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011101";
				elsif cntr ="001010011101" THEN
				      t1addb <= "00011101";
				      t2addb <= "00111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
						
				      
				      
				      
				      
				      
				      cntr <= "001010011110";
				elsif cntr ="001010011110" THEN
				      t1addb <= "00011110";
				      t2addb <= "00111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011111";
				elsif cntr ="001010011111" THEN
				      t1addb <= "00011111";
				      t2addb <= "00111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100000";
				elsif cntr ="001010100000" THEN
				      t1addb <= "00100000";
				      t2addb <= "00000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100001";
				elsif cntr ="001010100001" THEN
				      t1addb <= "00100001";
				      t2addb <= "00000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100010";
				elsif cntr ="001010100010" THEN
				      t1addb <= "00100010";
				      t2addb <= "00000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100011";
				elsif cntr ="001010100011" THEN
				      t1addb <= "00100011";
				      t2addb <= "00000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100100";
				elsif cntr ="001010100100" THEN
				      t1addb <= "00100100";		
				      t2addb <= "00000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100101";
				elsif cntr ="001010100101" THEN
				      t1addb <= "00100101";
				      t2addb <= "00000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100110";
				elsif cntr ="001010100110" THEN
				      t1addb <= "00100110";
				      t2addb <= "00000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100111";
				elsif cntr ="001010100111" THEN
				      t1addb <= "00100111";
				      t2addb <= "00000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101000";
				elsif cntr ="001010101000" THEN
				      t1addb <= "00101000";
				      t2addb <= "00001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101001";
				elsif cntr ="001010101001" THEN
				      t1addb <= "00101001";
				      t2addb <= "00001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101010";
				elsif cntr ="001010101010" THEN
				      t1addb <= "00101010";
				      t2addb <= "00001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
						
				      
				      cntr <= "001010101011";
				elsif cntr ="001010101011" THEN
				      t1addb <= "00101011";
				      t2addb <= "00001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101100";
				elsif cntr ="001010101100" THEN
				      t1addb <= "00101100";
				      t2addb <= "00001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101101";
				elsif cntr ="001010101101" THEN
				      t1addb <= "00101101";
				      t2addb <= "00001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101110";
				elsif cntr ="001010101110" THEN
				      t1addb <= "00101110";
				      t2addb <= "00001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;		
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101111";
				elsif cntr ="001010101111" THEN
				      t1addb <= "00101111";
				      t2addb <= "00001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110000";
				elsif cntr ="001010110000" THEN
				      t1addb <= "00110000";
				      t2addb <= "00010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110001";
				elsif cntr ="001010110001" THEN
				      t1addb <= "00110001";
				      t2addb <= "00010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110010";
				elsif cntr ="001010110010" THEN
				      t1addb <= "00110010";
				      t2addb <= "00010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110011";
				elsif cntr ="001010110011" THEN
				      t1addb <= "00110011";
				      t2addb <= "00010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110100";
				elsif cntr ="001010110100" THEN
				      t1addb <= "00110100";
				      t2addb <= "00010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110101";
				elsif cntr ="001010110101" THEN		
				      t1addb <= "00110101";
				      t2addb <= "00010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110110";
				elsif cntr ="001010110110" THEN
				      t1addb <= "00110110";
				      t2addb <= "00010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110111";
				elsif cntr ="001010110111" THEN
				      t1addb <= "00110111";
				      t2addb <= "00010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111000";
				elsif cntr ="001010111000" THEN
				      t1addb <= "00111000";
				      t2addb <= "00011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
						
				      
				      
				      
				      cntr <= "001010111001";
				elsif cntr ="001010111001" THEN
				      t1addb <= "00111001";
				      t2addb <= "00011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111010";
				elsif cntr ="001010111010" THEN
				      t1addb <= "00111010";
				      t2addb <= "00011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111011";
				elsif cntr ="001010111011" THEN
				      t1addb <= "00111011";
				      t2addb <= "00011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
						
				      
				      
				      cntr <= "001010111100";
				elsif cntr ="001010111100" THEN
				      t1addb <= "00111100";
				      t2addb <= "00011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111101";
				elsif cntr ="001010111101" THEN
				      t1addb <= "00111101";
				      t2addb <= "00011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111110";
				elsif cntr ="001010111110" THEN
				      t1addb <= "00111110";
				      t2addb <= "00011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111111";
				elsif cntr ="001010111111" THEN
				      t1addb <= "00111111";
				      t2addb <= "00011111";
				      bfrjin     <= t2doutb;		
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000000";
				elsif cntr ="001011000000" THEN
				      t1addb <= "01000000";
				      t2addb <= "01100000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000001";
				elsif cntr ="001011000001" THEN
				      t1addb <= "01000001";
				      t2addb <= "01100001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000010";
				      cntr <= "001011000010";
				elsif cntr ="001011000010" THEN
				      t1addb <= "01000010";
				      t2addb <= "01100010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000011";
				elsif cntr ="001011000011" THEN
				      t1addb <= "01000011";
				      t2addb <= "01100011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000100";
				elsif cntr ="001011000100" THEN
				      t1addb <= "01000100";
				      t2addb <= "01100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000101";
				elsif cntr ="001011000101" THEN
				      t1addb <= "01000101";
				      t2addb <= "01100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000110";		
				elsif cntr ="001011000110" THEN
				      t1addb <= "01000110";
				      t2addb <= "01100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000111";
				elsif cntr ="001011000111" THEN
				      t1addb <= "01000111";
				      t2addb <= "01100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001000";
				elsif cntr ="001011001000" THEN
				      t1addb <= "01001000";
				      t2addb <= "01101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001001";
				elsif cntr ="001011001001" THEN
				      t1addb <= "01001001";
				      t2addb <= "01101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
						
				      
				      
				      
				      
				      cntr <= "001011001010";
				elsif cntr ="001011001010" THEN
				      t1addb <= "01001010";
				      t2addb <= "01101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001011";
				elsif cntr ="001011001011" THEN
				      t1addb <= "01001011";
				      t2addb <= "01101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001100";
				elsif cntr ="001011001100" THEN
				      t1addb <= "01001100";
				      t2addb <= "01101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001101";
				elsif cntr ="001011001101" THEN
				      t1addb <= "01001101";
				      t2addb <= "01101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001110";
				elsif cntr ="001011001110" THEN
				      t1addb <= "01001110";
				      t2addb <= "01101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001111";
				elsif cntr ="001011001111" THEN
				      t1addb <= "01001111";
				      t2addb <= "01101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010000";
				elsif cntr ="001011010000" THEN
				      t1addb <= "01010000";
				      t2addb <= "01110000";		
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010001";
				elsif cntr ="001011010001" THEN
				      t1addb <= "01010001";
				      t2addb <= "01110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010010";
				elsif cntr ="001011010010" THEN
				      t1addb <= "01010010";
				      t2addb <= "01110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010011";
				elsif cntr ="001011010011" THEN
				      t1addb <= "01010011";
				      t2addb <= "01110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010100";
				elsif cntr ="001011010100" THEN
				      t1addb <= "01010100";
				      t2addb <= "01110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010101";
				elsif cntr ="001011010101" THEN
				      t1addb <= "01010101";
				      t2addb <= "01110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010110";
				elsif cntr ="001011010110" THEN
				      t1addb <= "01010110";
				      t2addb <= "01110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
						
				      cntr <= "001011010111";
				elsif cntr ="001011010111" THEN
				      t1addb <= "01010111";
				      t2addb <= "01110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011000";
				elsif cntr ="001011011000" THEN
				      t1addb <= "01011000";
				      t2addb <= "01111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011001";
				elsif cntr ="001011011001" THEN
				      t1addb <= "01011001";
				      t2addb <= "01111001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011010";
				elsif cntr ="001011011010" THEN
				      t1addb <= "01011010";
				      t2addb <= "01111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
						
				      
				      
				      
				      
				      
				      cntr <= "001011011011";
				elsif cntr ="001011011011" THEN
				      t1addb <= "01011011";
				      t2addb <= "01111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011100";
				elsif cntr ="001011011100" THEN
				      t1addb <= "01011100";
				      t2addb <= "01111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011101";
				elsif cntr ="001011011101" THEN
				      t1addb <= "01011101";
				      t2addb <= "01111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011110";
				elsif cntr ="001011011110" THEN
				      t1addb <= "01011110";
				      t2addb <= "01111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011111";
				elsif cntr ="001011011111" THEN
				      t1addb <= "01011111";
				      t2addb <= "01111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100000";
				elsif cntr ="001011100000" THEN
				      t1addb <= "01100000";
				      t2addb <= "01000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100001";
				elsif cntr ="001011100001" THEN
				      t1addb <= "01100001";		
				      t2addb <= "01000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100010";
				elsif cntr ="001011100010" THEN
				      t1addb <= "01100010";
				      t2addb <= "01000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100011";
				elsif cntr ="001011100011" THEN
				      t1addb <= "01100011";
				      t2addb <= "01000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100100";
				elsif cntr ="001011100100" THEN
				      t1addb <= "01100100";
				      t2addb <= "01000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100101";
				elsif cntr ="001011100101" THEN
				      t1addb <= "01100101";
				      t2addb <= "01000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100110";
				elsif cntr ="001011100110" THEN
				      t1addb <= "01100110";
				      t2addb <= "01000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100111";
				elsif cntr ="001011100111" THEN
				      t1addb <= "01100111";
				      t2addb <= "01000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
						
				      
				      cntr <= "001011101000";
				elsif cntr ="001011101000" THEN
				      t1addb <= "01101000";
				      t2addb <= "01001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101001";
				elsif cntr ="001011101001" THEN
				      t1addb <= "01101001";
				      t2addb <= "01001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101010";
				elsif cntr ="001011101010" THEN
				      t1addb <= "01101010";
				      t2addb <= "01001010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101011";
				elsif cntr ="001011101011" THEN
				      t1addb <= "01101011";
				      t2addb <= "01001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;		
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101100";
				elsif cntr ="001011101100" THEN
				      t1addb <= "01101100";
				      t2addb <= "01001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101101";
				elsif cntr ="001011101101" THEN
				      t1addb <= "01101101";
				      t2addb <= "01001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101110";
				elsif cntr ="001011101110" THEN
				      t1addb <= "01101110";
				      t2addb <= "01001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101111";
				elsif cntr ="001011101111" THEN
				      t1addb <= "01101111";
				      t2addb <= "01001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110000";
				elsif cntr ="001011110000" THEN
				      t1addb <= "01110000";
				      t2addb <= "01010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110001";
				elsif cntr ="001011110001" THEN
				      t1addb <= "01110001";
				      t2addb <= "01010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110010";
				elsif cntr ="001011110010" THEN		
				      t1addb <= "01110010";
				      t2addb <= "01010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110011";
				elsif cntr ="001011110011" THEN
				      t1addb <= "01110011";
				      t2addb <= "01010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110100";
				elsif cntr ="001011110100" THEN
				      t1addb <= "01110100";
				      t2addb <= "01010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110101";
				elsif cntr ="001011110101" THEN
				      t1addb <= "01110101";
				      t2addb <= "01010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
						
				      
				      
				      
				      cntr <= "001011110110";
				elsif cntr ="001011110110" THEN
				      t1addb <= "01110110";
				      t2addb <= "01010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110111";
				elsif cntr ="001011110111" THEN
				      t1addb <= "01110111";
				      t2addb <= "01010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111000";
				elsif cntr ="001011111000" THEN
				      t1addb <= "01111000";
				      t2addb <= "01011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
						
				      
				      
				      cntr <= "001011111001";
				elsif cntr ="001011111001" THEN
				      t1addb <= "01111001";
				      t2addb <= "01011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111010";
				elsif cntr ="001011111010" THEN
				      t1addb <= "01111010";
				      t2addb <= "01011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111011";
				elsif cntr ="001011111011" THEN
				      t1addb <= "01111011";
				      t2addb <= "01011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111100";
				elsif cntr ="001011111100" THEN
				      t1addb <= "01111100";
				      t2addb <= "01011100";
				      bfrjin     <= t2doutb;		
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111101";
				elsif cntr ="001011111101" THEN
				      t1addb <= "01111101";
				      t2addb <= "01011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111110";
				elsif cntr ="001011111110" THEN
				      t1addb <= "01111110";
				      t2addb <= "01011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111111";
				elsif cntr ="001011111111" THEN
				      t1addb <= "01111111";
				      t2addb <= "01011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000000";
				elsif cntr ="001100000000" THEN												
				      t1addb <= "10000000";      
				      t2addb <= "11000000";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000001";
				elsif cntr ="001100000001" THEN				
				      t1addb <= "10000001";      
				      t2addb <= "11000001";      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				        zetain   <="00000000";      
				      cntr <= "001100000010";
				elsif cntr ="001100000010" THEN		
				      t1addb <= "10000010";      
				      t2addb <= "11000010";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "001100000011";		
				elsif cntr ="001100000011" THEN		      
				      t1addb <= "10000011";      
				      t2addb <= "11000011";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001100000100";		      
				elsif cntr ="001100000100" THEN		       
				      t1addb <= "10000100";      
				      t2addb <= "11000100";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001100000101";	      
				elsif cntr ="001100000101" THEN	      
				      t1addb <= "10000101";      
				      t2addb <= "11000101";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001100000110";	           
				elsif cntr ="001100000110" THEN	           
				      t1addb <= "10000110";      
				      t2addb <= "11000110";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
						
				      
				                                    
				                                    
				                                    
				       cntr <= "001100000111";	      
				 elsif cntr ="001100000111" THEN	      
				      t1addb <= "10000111";      
				      t2addb <= "11000111";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                          
				                                          
				                                          
				       cntr <= "001100001000";	          
				 elsif cntr ="001100001000" THEN	      
				      t1addb <= "10001000";      
				      t2addb <= "11001000";      
				      bfrjin     <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				                                          
				                                          
				                                          
				      cntr <= "001100001001";	           										
				elsif cntr ="001100001001" THEN	 
				      t1addb <= "10001001";
				      t2addb <= "11001001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "001100001010";
				elsif cntr ="001100001010" THEN
				      t1addb <= "10001010";
				      t2addb <= "11001010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001011";
				elsif cntr ="001100001011" THEN
				      t1addb <= "10001011";
				      t2addb <= "11001011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001100";
				elsif cntr ="001100001100" THEN
				      t1addb <= "10001100";
				      t2addb <= "11001100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001101";
				elsif cntr ="001100001101" THEN
				      t1addb <= "10001101";
				      t2addb <= "11001101";		
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001110";
				elsif cntr ="001100001110" THEN
				      t1addb <= "10001110";
				      t2addb <= "11001110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001111";
				elsif cntr ="001100001111" THEN
				      t1addb <= "10001111";
				      t2addb <= "11001111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010000";
				elsif cntr ="001100010000" THEN
				      t1addb <= "10010000";
				      t2addb <= "11010000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010001";
				elsif cntr ="001100010001" THEN
				      t1addb <= "10010001";
				      t2addb <= "11010001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010010";
				elsif cntr ="001100010010" THEN
				      t1addb <= "10010010";
				      t2addb <= "11010010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010011";
				elsif cntr ="001100010011" THEN
				      t1addb <= "10010011";
				      t2addb <= "11010011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
						
				      cntr <= "001100010100";
				elsif cntr ="001100010100" THEN
				      t1addb <= "10010100";
				      t2addb <= "11010100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010101";
				elsif cntr ="001100010101" THEN
				      t1addb <= "10010101";
				      t2addb <= "11010101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010110";
				elsif cntr ="001100010110" THEN
				      t1addb <= "10010110";
				      t2addb <= "11010110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010111";
				elsif cntr ="001100010111" THEN
				      t1addb <= "10010111";
				      t2addb <= "11010111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
						
				      
				      
				      
				      
				      
				      cntr <= "001100011000";
				elsif cntr ="001100011000" THEN
				      t1addb <= "10011000";
				      t2addb <= "11011000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011001";
				elsif cntr ="001100011001" THEN
				      t1addb <= "10011001";
				      t2addb <= "11011001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011010";
				elsif cntr ="001100011010" THEN
				      t1addb <= "10011010";
				      t2addb <= "11011010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011011";
				elsif cntr ="001100011011" THEN
				      t1addb <= "10011011";
				      t2addb <= "11011011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011100";
				elsif cntr ="001100011100" THEN
				      t1addb <= "10011100";
				      t2addb <= "11011100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011101";
				elsif cntr ="001100011101" THEN
				      t1addb <= "10011101";
				      t2addb <= "11011101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011110";
				elsif cntr ="001100011110" THEN
				      t1addb <= "10011110";		
				      t2addb <= "11011110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011111";
				elsif cntr ="001100011111" THEN
				      t1addb <= "10011111";
				      t2addb <= "11011111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100000";
				elsif cntr ="001100100000" THEN
				      t1addb <= "10100000";
				      t2addb <= "11100000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100001";
				elsif cntr ="001100100001" THEN
				      t1addb <= "10100001";
				      t2addb <= "11100001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100010";
				elsif cntr ="001100100010" THEN
				      t1addb <= "10100010";
				      t2addb <= "11100010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100011";
				elsif cntr ="001100100011" THEN
				      t1addb <= "10100011";
				      t2addb <= "11100011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100100";
				elsif cntr ="001100100100" THEN
				      t1addb <= "10100100";
				      t2addb <= "11100100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
						
				      
				      cntr <= "001100100101";
				elsif cntr ="001100100101" THEN
				      t1addb <= "10100101";
				      t2addb <= "11100101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100110";
				elsif cntr ="001100100110" THEN
				      t1addb <= "10100110";
				      t2addb <= "11100110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100111";
				elsif cntr ="001100100111" THEN
				      t1addb <= "10100111";
				      t2addb <= "11100111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101000";
				elsif cntr ="001100101000" THEN
				      t1addb <= "10101000";
				      t2addb <= "11101000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;		
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101001";
				elsif cntr ="001100101001" THEN
				      t1addb <= "10101001";
				      t2addb <= "11101001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101010";
				elsif cntr ="001100101010" THEN
				      t1addb <= "10101010";
				      t2addb <= "11101010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101011";
				elsif cntr ="001100101011" THEN
				      t1addb <= "10101011";
				      t2addb <= "11101011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101100";
				elsif cntr ="001100101100" THEN
				      t1addb <= "10101100";
				      t2addb <= "11101100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101101";
				elsif cntr ="001100101101" THEN
				      t1addb <= "10101101";
				      t2addb <= "11101101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101110";
				elsif cntr ="001100101110" THEN
				      t1addb <= "10101110";
				      t2addb <= "11101110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101111";
				elsif cntr ="001100101111" THEN		
				      t1addb <= "10101111";
				      t2addb <= "11101111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110000";
				elsif cntr ="001100110000" THEN
				      t1addb <= "10110000";
				      t2addb <= "11110000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110001";
				elsif cntr ="001100110001" THEN
				      t1addb <= "10110001";
				      t2addb <= "11110001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110010";
				elsif cntr ="001100110010" THEN
				      t1addb <= "10110010";
				      t2addb <= "11110010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
						
				      
				      
				      
				      cntr <= "001100110011";
				elsif cntr ="001100110011" THEN
				      t1addb <= "10110011";
				      t2addb <= "11110011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110100";
				elsif cntr ="001100110100" THEN
				      t1addb <= "10110100";
				      t2addb <= "11110100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110101";
				elsif cntr ="001100110101" THEN
				      t1addb <= "10110101";
				      t2addb <= "11110101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
						
				      
				      
				      cntr <= "001100110110";
				elsif cntr ="001100110110" THEN
				      t1addb <= "10110110";
				      t2addb <= "11110110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110111";
				elsif cntr ="001100110111" THEN
				      t1addb <= "10110111";
				      t2addb <= "11110111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111000";
				elsif cntr ="001100111000" THEN
				      t1addb <= "10111000";
				      t2addb <= "11111000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111001";
				elsif cntr ="001100111001" THEN
				      t1addb <= "10111001";
				      t2addb <= "11111001";
				      bfrjin     <= t1doutb;		
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111010";
				elsif cntr ="001100111010" THEN
				      t1addb <= "10111010";
				      t2addb <= "11111010";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111011";
				elsif cntr ="001100111011" THEN
				      t1addb <= "10111011";
				      t2addb <= "11111011";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111100";
				elsif cntr ="001100111100" THEN
				      t1addb <= "10111100";
				      t2addb <= "11111100";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111101";
				elsif cntr ="001100111101" THEN
				      t1addb <= "10111101";
				      t2addb <= "11111101";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111110";
				elsif cntr ="001100111110" THEN
				      t1addb <= "10111110";
				      t2addb <= "11111110";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111111";
				elsif cntr ="001100111111" THEN
				      t1addb <= "10111111";
				      t2addb <= "11111111";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000000";		
				elsif cntr ="001101000000" THEN
				      t1addb <= "11000000";
				      t2addb <= "10000000";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000001";
				elsif cntr ="001101000001" THEN
				      t1addb <= "11000001";
				      t2addb <= "10000001";
				      bfrjin     <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000010";
				elsif cntr ="001101000010" THEN
				      t1addb <= "11000010";
				      t2addb <= "10000010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000011";
				elsif cntr ="001101000011" THEN
				      t1addb <= "11000011";
				      t2addb <= "10000011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
						
				      
				      
				      
				      
				      cntr <= "001101000100";
				elsif cntr ="001101000100" THEN
				      t1addb <= "11000100";
				      t2addb <= "10000100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000101";
				elsif cntr ="001101000101" THEN
				      t1addb <= "11000101";
				      t2addb <= "10000101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000110";
				elsif cntr ="001101000110" THEN
				      t1addb <= "11000110";
				      t2addb <= "10000110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000111";
				elsif cntr ="001101000111" THEN
				      t1addb <= "11000111";
				      t2addb <= "10000111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001000";
				elsif cntr ="001101001000" THEN
				      t1addb <= "11001000";
				      t2addb <= "10001000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001001";
				elsif cntr ="001101001001" THEN
				      t1addb <= "11001001";
				      t2addb <= "10001001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001010";
				elsif cntr ="001101001010" THEN
				      t1addb <= "11001010";
				      t2addb <= "10001010";		
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001011";
				elsif cntr ="001101001011" THEN
				      t1addb <= "11001011";
				      t2addb <= "10001011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001100";
				elsif cntr ="001101001100" THEN
				      t1addb <= "11001100";
				      t2addb <= "10001100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001101";
				elsif cntr ="001101001101" THEN
				      t1addb <= "11001101";
				      t2addb <= "10001101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001110";
				elsif cntr ="001101001110" THEN
				      t1addb <= "11001110";
				      t2addb <= "10001110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001111";
				elsif cntr ="001101001111" THEN
				      t1addb <= "11001111";
				      t2addb <= "10001111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010000";
				elsif cntr ="001101010000" THEN
				      t1addb <= "11010000";
				      t2addb <= "10010000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
						
				      cntr <= "001101010001";
				elsif cntr ="001101010001" THEN
				      t1addb <= "11010001";
				      t2addb <= "10010001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010010";
				elsif cntr ="001101010010" THEN
				      t1addb <= "11010010";
				      t2addb <= "10010010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010011";
				elsif cntr ="001101010011" THEN
				      t1addb <= "11010011";
				      t2addb <= "10010011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010100";
				elsif cntr ="001101010100" THEN
				      t1addb <= "11010100";
				      t2addb <= "10010100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
						
				      
				      
				      
				      
				      
				      cntr <= "001101010101";
				elsif cntr ="001101010101" THEN
				      t1addb <= "11010101";
				      t2addb <= "10010101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010110";
				elsif cntr ="001101010110" THEN
				      t1addb <= "11010110";
				      t2addb <= "10010110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010111";
				elsif cntr ="001101010111" THEN
				      t1addb <= "11010111";
				      t2addb <= "10010111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011000";
				elsif cntr ="001101011000" THEN
				      t1addb <= "11011000";
				      t2addb <= "10011000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011001";
				elsif cntr ="001101011001" THEN
				      t1addb <= "11011001";
				      t2addb <= "10011001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011010";
				elsif cntr ="001101011010" THEN
				      t1addb <= "11011010";
				      t2addb <= "10011010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011011";
				elsif cntr ="001101011011" THEN
				      t1addb <= "11011011";		
				      t2addb <= "10011011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011100";
				elsif cntr ="001101011100" THEN
				      t1addb <= "11011100";
				      t2addb <= "10011100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011101";
				elsif cntr ="001101011101" THEN
				      t1addb <= "11011101";
				      t2addb <= "10011101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011110";
				elsif cntr ="001101011110" THEN
				      t1addb <= "11011110";
				      t2addb <= "10011110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011111";
				elsif cntr ="001101011111" THEN
				      t1addb <= "11011111";
				      t2addb <= "10011111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100000";
				elsif cntr ="001101100000" THEN
				      t1addb <= "11100000";
				      t2addb <= "10100000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100001";
				elsif cntr ="001101100001" THEN
				      t1addb <= "11100001";
				      t2addb <= "10100001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
						
				      
				      cntr <= "001101100010";
				elsif cntr ="001101100010" THEN
				      t1addb <= "11100010";
				      t2addb <= "10100010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100011";
				elsif cntr ="001101100011" THEN
				      t1addb <= "11100011";
				      t2addb <= "10100011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100100";
				elsif cntr ="001101100100" THEN
				      t1addb <= "11100100";
				      t2addb <= "10100100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100101";
				elsif cntr ="001101100101" THEN
				      t1addb <= "11100101";
				      t2addb <= "10100101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;		
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100110";
				elsif cntr ="001101100110" THEN
				      t1addb <= "11100110";
				      t2addb <= "10100110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100111";
				elsif cntr ="001101100111" THEN
				      t1addb <= "11100111";
				      t2addb <= "10100111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101000";
				elsif cntr ="001101101000" THEN
				      t1addb <= "11101000";
				      t2addb <= "10101000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101001";
				elsif cntr ="001101101001" THEN
				      t1addb <= "11101001";
				      t2addb <= "10101001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101010";
				elsif cntr ="001101101010" THEN
				      t1addb <= "11101010";
				      t2addb <= "10101010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101011";
				elsif cntr ="001101101011" THEN
				      t1addb <= "11101011";
				      t2addb <= "10101011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101100";
				elsif cntr ="001101101100" THEN		
				      t1addb <= "11101100";
				      t2addb <= "10101100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101101";
				elsif cntr ="001101101101" THEN
				      t1addb <= "11101101";
				      t2addb <= "10101101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101110";
				elsif cntr ="001101101110" THEN
				      t1addb <= "11101110";
				      t2addb <= "10101110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101111";
				elsif cntr ="001101101111" THEN
				      t1addb <= "11101111";
				      t2addb <= "10101111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
						
				      
				      
				      
				      cntr <= "001101110000";
				elsif cntr ="001101110000" THEN
				      t1addb <= "11110000";
				      t2addb <= "10110000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110001";
				elsif cntr ="001101110001" THEN
				      t1addb <= "11110001";
				      t2addb <= "10110001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110010";
				elsif cntr ="001101110010" THEN
				      t1addb <= "11110010";
				      t2addb <= "10110010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
						
				      
				      
				      cntr <= "001101110011";
				elsif cntr ="001101110011" THEN
				      t1addb <= "11110011";
				      t2addb <= "10110011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110100";
				elsif cntr ="001101110100" THEN
				      t1addb <= "11110100";
				      t2addb <= "10110100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110101";
				elsif cntr ="001101110101" THEN
				      t1addb <= "11110101";
				      t2addb <= "10110101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110110";
				elsif cntr ="001101110110" THEN
				      t1addb <= "11110110";
				      t2addb <= "10110110";
				      bfrjin     <= t2doutb;		
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110111";
				elsif cntr ="001101110111" THEN
				      t1addb <= "11110111";
				      t2addb <= "10110111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111000";
				elsif cntr ="001101111000" THEN
				      t1addb <= "11111000";
				      t2addb <= "10111000";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111001";
				elsif cntr ="001101111001" THEN
				      t1addb <= "11111001";
				      t2addb <= "10111001";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111010";
				elsif cntr ="001101111010" THEN
				      t1addb <= "11111010";
				      t2addb <= "10111010";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111011";
				elsif cntr ="001101111011" THEN
				      t1addb <= "11111011";
				      t2addb <= "10111011";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111100";
				elsif cntr ="001101111100" THEN
				      t1addb <= "11111100";
				      t2addb <= "10111100";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111101";		
				elsif cntr ="001101111101" THEN
				      t1addb <= "11111101";
				      t2addb <= "10111101";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111110";
				elsif cntr ="001101111110" THEN
				      t1addb <= "11111110";
				      t2addb <= "10111110";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111111";
				elsif cntr ="001101111111" THEN
				      t1addb <= "11111111";
				      t2addb <= "10111111";
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000000";
				elsif cntr ="001110000000" THEN												
				      t1addb <= "00000000";      
				      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
						
				      
				      
				      
				      
				      cntr <= "001110000001";
				elsif cntr ="001110000001" THEN	
				      t1addb <= "00000001";      
				      
				      bfrjin     <= t2doutb;
				      bfrjplin <= t1doutb;
				      
						
				      
				      
				      
				        zetain   <="10000000";      
				      cntr <= "001110000010";
				elsif cntr ="001110000010" THEN	
				      t1addb <= "00000010";      
				      
				      bfrjplin     <= t1doutb;      
				      bfrjin <= "000000000000";
				      
				      
				      
				            
				            
				            
				      cntr <= "001110000011";      
				elsif cntr ="001110000011" THEN	      
				      t1addb <= "00000011";      
				      
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001110000100";           
				elsif cntr ="001110000100" THEN	        
				      t1addb <= "00000100";      
				      
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001110000101";             
				elsif cntr ="001110000101" THEN	          
				      t1addb <= "00000101";      
				      
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001110000110";                
				elsif cntr ="001110000110" THEN	             
				      t1addb <= "00000110";      
				      
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001110000111";            
				elsif cntr ="001110000111" THEN	         
				      t1addb <= "00000111";      
						
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                                          
				                                          
				                                          
				      cntr <= "001110001000";                  
				elsif cntr ="001110001000" THEN	               
				      t1addb <= "00001000";      
				      
				      bfrjplin     <= t1doutb;      
				      
				      
				      
				      
				                                   
				                                   
				                                   
				      cntr <= "001110001001";      
				elsif cntr ="001110001001" THEN	   
				      t1addb <= "00001001";
				
				      bfrjplin     <= t1doutb;
				
					  
				
				
					  
				      
				      
				      
				      cntr <= "001110001010";
				elsif cntr ="001110001010" THEN
				      t1addb <= "00001010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001011";
				elsif cntr ="001110001011" THEN
				      t1addb <= "00001011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001100";
				elsif cntr ="001110001100" THEN
				      t1addb <= "00001100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001101";
				elsif cntr ="001110001101" THEN
				      t1addb <= "00001101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
						
				      cntr <= "001110001110";
				elsif cntr ="001110001110" THEN
				      t1addb <= "00001110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001111";
				elsif cntr ="001110001111" THEN
				      t1addb <= "00001111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010000";
				elsif cntr ="001110010000" THEN
				      t1addb <= "00010000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010001";
				elsif cntr ="001110010001" THEN
				      t1addb <= "00010001";
				      
				      bfrjplin     <= t1doutb;
				      
						
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010010";
				elsif cntr ="001110010010" THEN
				      t1addb <= "00010010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010011";
				elsif cntr ="001110010011" THEN
				      t1addb <= "00010011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010100";
				elsif cntr ="001110010100" THEN
				      t1addb <= "00010100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010101";
				elsif cntr ="001110010101" THEN
				      t1addb <= "00010101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010110";
				elsif cntr ="001110010110" THEN
				      t1addb <= "00010110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110010111";
				elsif cntr ="001110010111" THEN
				      t1addb <= "00010111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011000";
				elsif cntr ="001110011000" THEN
				      t1addb <= "00011000";		
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011001";
				elsif cntr ="001110011001" THEN
				      t1addb <= "00011001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011010";
				elsif cntr ="001110011010" THEN
				      t1addb <= "00011010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011011";
				elsif cntr ="001110011011" THEN
				      t1addb <= "00011011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
						
				      
				      
				      
				      cntr <= "001110011100";
				elsif cntr ="001110011100" THEN
				      t1addb <= "00011100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011101";
				elsif cntr ="001110011101" THEN
				      t1addb <= "00011101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110011110";
				elsif cntr ="001110011110" THEN
				      t1addb <= "00011110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
						
				      
				      cntr <= "001110011111";
				elsif cntr ="001110011111" THEN
				      t1addb <= "00011111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100000";
				elsif cntr ="001110100000" THEN
				      t1addb <= "00100000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100001";
				elsif cntr ="001110100001" THEN
				      t1addb <= "00100001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100010";
				elsif cntr ="001110100010" THEN
				      t1addb <= "00100010";
				      
				      bfrjplin     <= t1doutb;
						
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100011";
				elsif cntr ="001110100011" THEN
				      t1addb <= "00100011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100100";
				elsif cntr ="001110100100" THEN
				      t1addb <= "00100100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100101";
				elsif cntr ="001110100101" THEN
				      t1addb <= "00100101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100110";
				elsif cntr ="001110100110" THEN
				      t1addb <= "00100110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110100111";
				elsif cntr ="001110100111" THEN
				      t1addb <= "00100111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101000";
				elsif cntr ="001110101000" THEN
				      t1addb <= "00101000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101001";
				elsif cntr ="001110101001" THEN		
				      t1addb <= "00101001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101010";
				elsif cntr ="001110101010" THEN
				      t1addb <= "00101010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101011";
				elsif cntr ="001110101011" THEN
				      t1addb <= "00101011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101100";
				elsif cntr ="001110101100" THEN
				      t1addb <= "00101100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
						
				      
				      
				      
				      
				      cntr <= "001110101101";
				elsif cntr ="001110101101" THEN
				      t1addb <= "00101101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101110";
				elsif cntr ="001110101110" THEN
				      t1addb <= "00101110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110101111";
				elsif cntr ="001110101111" THEN
				      t1addb <= "00101111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
						
				      
				      
				      cntr <= "001110110000";
				elsif cntr ="001110110000" THEN
				      t1addb <= "00110000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110001";
				elsif cntr ="001110110001" THEN
				      t1addb <= "00110001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110010";
				elsif cntr ="001110110010" THEN
				      t1addb <= "00110010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110011";
				elsif cntr ="001110110011" THEN
				      t1addb <= "00110011";
				      
				      bfrjplin     <= t1doutb;		
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110100";
				elsif cntr ="001110110100" THEN
				      t1addb <= "00110100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110101";
				elsif cntr ="001110110101" THEN
				      t1addb <= "00110101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110110";
				elsif cntr ="001110110110" THEN
				      t1addb <= "00110110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110110111";
				elsif cntr ="001110110111" THEN
				      t1addb <= "00110111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111000";
				elsif cntr ="001110111000" THEN
				      t1addb <= "00111000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111001";
				elsif cntr ="001110111001" THEN
				      t1addb <= "00111001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111010";		
				elsif cntr ="001110111010" THEN
				      t1addb <= "00111010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111011";
				elsif cntr ="001110111011" THEN
				      t1addb <= "00111011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111100";
				elsif cntr ="001110111100" THEN
				      t1addb <= "00111100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111101";
				elsif cntr ="001110111101" THEN
				      t1addb <= "00111101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
						
				      
				      
				      
				      
				      
				      cntr <= "001110111110";
				elsif cntr ="001110111110" THEN
				      t1addb <= "00111110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110111111";
				elsif cntr ="001110111111" THEN
				      t1addb <= "00111111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000000";
				elsif cntr ="001111000000" THEN
				      t1addb <= "01000000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000001";
				elsif cntr ="001111000001" THEN
				      t1addb <= "01000001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000010";
				elsif cntr ="001111000010" THEN
				      t1addb <= "01000010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000011";
				elsif cntr ="001111000011" THEN
				      t1addb <= "01000011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000100";
				elsif cntr ="001111000100" THEN
				      t1addb <= "01000100";
						
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000101";
				elsif cntr ="001111000101" THEN
				      t1addb <= "01000101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000110";
				elsif cntr ="001111000110" THEN
				      t1addb <= "01000110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111000111";
				elsif cntr ="001111000111" THEN
				      t1addb <= "01000111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001000";
				elsif cntr ="001111001000" THEN
				      t1addb <= "01001000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001001";
				elsif cntr ="001111001001" THEN
				      t1addb <= "01001001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001010";
				elsif cntr ="001111001010" THEN
				      t1addb <= "01001010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
						
				      cntr <= "001111001011";
				elsif cntr ="001111001011" THEN
				      t1addb <= "01001011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001100";
				elsif cntr ="001111001100" THEN
				      t1addb <= "01001100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001101";
				elsif cntr ="001111001101" THEN
				      t1addb <= "01001101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001110";
				elsif cntr ="001111001110" THEN
				      t1addb <= "01001110";
				      
				      bfrjplin     <= t1doutb;
				      
						
				      
				      
				      
				      
				      
				      
				      cntr <= "001111001111";
				elsif cntr ="001111001111" THEN
				      t1addb <= "01001111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010000";
				elsif cntr ="001111010000" THEN
				      t1addb <= "01010000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010001";
				elsif cntr ="001111010001" THEN
				      t1addb <= "01010001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010010";
				elsif cntr ="001111010010" THEN
				      t1addb <= "01010010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010011";
				elsif cntr ="001111010011" THEN
				      t1addb <= "01010011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010100";
				elsif cntr ="001111010100" THEN
				      t1addb <= "01010100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010101";
				elsif cntr ="001111010101" THEN
				      t1addb <= "01010101";		
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010110";
				elsif cntr ="001111010110" THEN
				      t1addb <= "01010110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111010111";
				elsif cntr ="001111010111" THEN
				      t1addb <= "01010111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011000";
				elsif cntr ="001111011000" THEN
				      t1addb <= "01011000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
						
				      
				      
				      
				      cntr <= "001111011001";
				elsif cntr ="001111011001" THEN
				      t1addb <= "01011001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011010";
				elsif cntr ="001111011010" THEN
				      t1addb <= "01011010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011011";
				elsif cntr ="001111011011" THEN
				      t1addb <= "01011011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
						
				      
				      cntr <= "001111011100";
				elsif cntr ="001111011100" THEN
				      t1addb <= "01011100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011101";
				elsif cntr ="001111011101" THEN
				      t1addb <= "01011101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011110";
				elsif cntr ="001111011110" THEN
				      t1addb <= "01011110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111011111";
				elsif cntr ="001111011111" THEN
				      t1addb <= "01011111";
				      
				      bfrjplin     <= t1doutb;
						
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100000";
				elsif cntr ="001111100000" THEN
				      t1addb <= "01100000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100001";
				elsif cntr ="001111100001" THEN
				      t1addb <= "01100001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100010";
				elsif cntr ="001111100010" THEN
				      t1addb <= "01100010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100011";
				elsif cntr ="001111100011" THEN
				      t1addb <= "01100011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100100";
				elsif cntr ="001111100100" THEN
				      t1addb <= "01100100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100101";
				elsif cntr ="001111100101" THEN
				      t1addb <= "01100101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100110";
				elsif cntr ="001111100110" THEN		
				      t1addb <= "01100110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111100111";
				elsif cntr ="001111100111" THEN
				      t1addb <= "01100111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101000";
				elsif cntr ="001111101000" THEN
				      t1addb <= "01101000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101001";
				elsif cntr ="001111101001" THEN
				      t1addb <= "01101001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
						
				      
				      
				      
				      
				      cntr <= "001111101010";
				elsif cntr ="001111101010" THEN
				      t1addb <= "01101010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101011";
				elsif cntr ="001111101011" THEN
				      t1addb <= "01101011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101100";
				elsif cntr ="001111101100" THEN
				      t1addb <= "01101100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
						
				      
				      
				      cntr <= "001111101101";
				elsif cntr ="001111101101" THEN
				      t1addb <= "01101101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101110";
				elsif cntr ="001111101110" THEN
				      t1addb <= "01101110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111101111";
				elsif cntr ="001111101111" THEN
				      t1addb <= "01101111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110000";
				elsif cntr ="001111110000" THEN
				      t1addb <= "01110000";
				      
				      bfrjplin     <= t1doutb;		
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110001";
				elsif cntr ="001111110001" THEN
				      t1addb <= "01110001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110010";
				elsif cntr ="001111110010" THEN
				      t1addb <= "01110010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110011";
				elsif cntr ="001111110011" THEN
				      t1addb <= "01110011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110100";
				elsif cntr ="001111110100" THEN
				      t1addb <= "01110100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110101";
				elsif cntr ="001111110101" THEN
				      t1addb <= "01110101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110110";
				elsif cntr ="001111110110" THEN
				      t1addb <= "01110110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111110111";		
				elsif cntr ="001111110111" THEN
				      t1addb <= "01110111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111000";
				elsif cntr ="001111111000" THEN
				      t1addb <= "01111000";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111001";
				elsif cntr ="001111111001" THEN
				      t1addb <= "01111001";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111010";
				elsif cntr ="001111111010" THEN
				      t1addb <= "01111010";
				      
				      bfrjplin     <= t1doutb;
				      
				      
						
				      
				      
				      
				      
				      
				      cntr <= "001111111011";
				elsif cntr ="001111111011" THEN
				      t1addb <= "01111011";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111100";
				elsif cntr ="001111111100" THEN
				      t1addb <= "01111100";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111101";
				elsif cntr ="001111111101" THEN
				      t1addb <= "01111101";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111110";
				elsif cntr ="001111111110" THEN
				      t1addb <= "01111110";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001111111111";
				elsif cntr ="001111111111" THEN
				      t1addb <= "01111111";
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "010000000000";
				elsif cntr ="010000000000" THEN
				      
				      
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "010000000001";
				elsif cntr ="010000000001" THEN
				      
						
				      bfrjplin     <= t1doutb;
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "010000000010";
				elsif cntr ="010000000010" THEN
				      
				      
				      
				      
				      
				      
				      
				      
				            
				            
				            
				      cntr <= "010000000011";      
				elsif cntr ="010000000011" THEN      
				      
				      
				      
				      
				      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "010000000100";           
				elsif cntr ="010000000100" THEN         
				      
				      
				      
				      
				      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "010000000101";          
				elsif cntr ="010000000101" THEN        
				      
				      
				      
				      
				      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "010000000110";            
				elsif cntr ="010000000110" THEN          
				      
				      
				      
				      
				      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "010000000111";          
				elsif cntr ="010000000111" THEN        
				      
				      
				      
				      
				      
				      
				      
				      
				                                        
				                                        
				                                  		
				      cntr <= "010000001000";           
				elsif cntr ="010000001000" THEN         
				      
				      
				      
				      
				      
				      
				      
				      
				                                    
				       
					
				                                  	
				      cntr <= "010000001001";       
				elsif cntr ="010000001001" THEN     
				
						
					 
				
				      cntr <= "010000001010";       
				elsif cntr ="010000001010" THEN 
				
					pdone <= '1';
				
				
				cntr <= "010000001011";       
				elsif cntr ="010000001011" THEN 
				
					  cntr <= "000000000000"; 
				
				
				
				
		
				
				END IF;





				
				IF cntr1 ="000000000000" THEN
					  
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000001" THEN
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000010" THEN
				
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000011" THEN
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000100" THEN
				
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000101" THEN
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000110" THEN
				
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000000111" THEN
				
				
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000001000" THEN
				
				
					  
				
				
				
				
				
				
				
				
				ELSIF cntr1 ="000000001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000000";
				      t2adda <= "00000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
				      t2adda <= "00000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
				      t2adda <= "00000010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
				      t2adda <= "00000011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000100";
				      t2adda <= "00000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
				      t2adda <= "00000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000111";
				      t2adda <= "00000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001000";
				      t2adda <= "00001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001010";
				      t2adda <= "00001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
				      t2adda <= "00001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
				      t2adda <= "00001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
				      t2adda <= "00001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001111";
				      t2adda <= "00001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010000";
				      t2adda <= "00010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010001";
				      t2adda <= "00010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010010";
				      t2adda <= "00010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010011";
				      t2adda <= "00010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010100";
				      t2adda <= "00010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010101";
				      t2adda <= "00010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010110";
				      t2adda <= "00010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010111";
				      t2adda <= "00010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011000";
				      t2adda <= "00011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
				      t2adda <= "00011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011100";
				      t2adda <= "00011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011101";
				      t2adda <= "00011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011110";
				      t2adda <= "00011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011111";
				      t2adda <= "00011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100000";
				      t2adda <= "00100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100001";
				      t2adda <= "00100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
				      t2adda <= "00100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100110";
				      t2adda <= "00100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100111";
				      t2adda <= "00100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101001";
				      t2adda <= "00101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101010";
				      t2adda <= "00101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101011";
				      t2adda <= "00101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101100";
				      t2adda <= "00101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101101";
				      t2adda <= "00101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101110";
				      t2adda <= "00101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101111";
				      t2adda <= "00101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110000";
				      t2adda <= "00110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110001";
				      t2adda <= "00110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
				      t2adda <= "00110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000000111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000000111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
				      t2adda <= "00110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000000111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
				      t2adda <= "00110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000000111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
				      t2adda <= "00110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111000";
				      t2adda <= "00111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
				      t2adda <= "00111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111010";
				      t2adda <= "00111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111011";
				      t2adda <= "00111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111100";
				      t2adda <= "00111100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111101";
				      t2adda <= "00111101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111110";
				      t2adda <= "00111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111111";
				      t2adda <= "00111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000000";
				      t2adda <= "01000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000001";
				      t2adda <= "01000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000010";
				      t2adda <= "01000010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000011";
				      t2adda <= "01000011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000100";
				      t2adda <= "01000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000101";
				      t2adda <= "01000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000110";
				      t2adda <= "01000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
				      t2adda <= "01000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001000";
				      t2adda <= "01001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
				      t2adda <= "01001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001010";
				      t2adda <= "01001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
				      t2adda <= "01001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001100";
				      t2adda <= "01001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001101";
				      t2adda <= "01001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001110";
				      t2adda <= "01001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001111";
				      t2adda <= "01001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010000";
				      t2adda <= "01010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010001";
				      t2adda <= "01010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
				      t2adda <= "01010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010011";
				      t2adda <= "01010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
				      t2adda <= "01010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
				      t2adda <= "01010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
				      t2adda <= "01010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
				      t2adda <= "01010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
				      t2adda <= "01011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011001";
				      t2adda <= "01011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
				      t2adda <= "01011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
				      t2adda <= "01011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
				      t2adda <= "01011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011101";
				      t2adda <= "01011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011110";
				      t2adda <= "01011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011111";
				      t2adda <= "01011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
				      t2adda <= "01100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100010";
				      t2adda <= "01100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100011";
				      t2adda <= "01100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100100";
				      t2adda <= "01100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100101";
				      t2adda <= "01100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100110";
				      t2adda <= "01100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100111";
				      t2adda <= "01100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
				      t2adda <= "01101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101001";
				      t2adda <= "01101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
				      t2adda <= "01101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
				      t2adda <= "01101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101101";
				      t2adda <= "01101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101110";
				      t2adda <= "01101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101111";
				      t2adda <= "01101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110000";
				      t2adda <= "01110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110001";
				      t2adda <= "01110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
				      t2adda <= "01110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000001111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110011";
				      t2adda <= "01110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000001111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110100";
				      t2adda <= "01110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000001111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110101";
				      t2adda <= "01110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				ELSIF cntr1 ="000001111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110110";
				      t2adda <= "01110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				ELSIF cntr1 ="000010000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110111";
				      t2adda <= "01110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				ELSIF cntr1 ="000010000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111000";
				      t2adda <= "01111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				ELSIF cntr1 ="000010000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111001";
				      t2adda <= "01111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				            
				            
				            
				ELSIF cntr1 ="000010000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111010";
				      t2adda <= "01111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				ELSIF cntr1 ="000010000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111011";
				      t2adda <= "01111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				ELSIF cntr1 ="000010000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111100";
				      t2adda <= "01111100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				                              
				                              
				ELSIF cntr1 ="000010000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111101";
				      t2adda <= "01111101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				                                    
				                                    
				                                    
				ELSIF cntr1 ="000010000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111110";
				      t2adda <= "01111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                          
				                                          
				                                          
				ELSIF cntr1 ="000010001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111111";
				      t2adda <= "01111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                         
				                                         										
				                                   
				ELSIF cntr1 ="000010001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000000";
				      t2adda <= "10000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000001";
				      t2adda <= "10000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000010";
				      t2adda <= "10000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000011";
				      t2adda <= "10000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000100";
				      t2adda <= "10000100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000101";
				      t2adda <= "10000101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000110";
				      t2adda <= "10000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000111";
				      t2adda <= "10000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001000";
				      t2adda <= "10001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001001";
				      t2adda <= "10001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001010";
				      t2adda <= "10001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001011";
				      t2adda <= "10001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001100";
				      t2adda <= "10001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001101";
				      t2adda <= "10001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001110";
				      t2adda <= "10001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001111";
				      t2adda <= "10001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010000";
				      t2adda <= "10010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010001";
				      t2adda <= "10010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010010";
				      t2adda <= "10010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010011";
				      t2adda <= "10010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010100";
				      t2adda <= "10010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010101";
				      t2adda <= "10010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010110";
				      t2adda <= "10010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010111";
				      t2adda <= "10010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011000";
				      t2adda <= "10011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011001";
				      t2adda <= "10011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011010";
				      t2adda <= "10011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011011";
				      t2adda <= "10011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011100";
				      t2adda <= "10011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011101";
				      t2adda <= "10011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011110";
				      t2adda <= "10011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011111";
				      t2adda <= "10011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100000";
				      t2adda <= "10100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100001";
				      t2adda <= "10100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100010";
				      t2adda <= "10100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100011";
				      t2adda <= "10100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100100";
				      t2adda <= "10100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100101";
				      t2adda <= "10100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100110";
				      t2adda <= "10100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100111";
				      t2adda <= "10100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101000";
				      t2adda <= "10101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101001";
				      t2adda <= "10101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101010";
				      t2adda <= "10101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101011";
				      t2adda <= "10101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101100";
				      t2adda <= "10101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101101";
				      t2adda <= "10101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101110";
				      t2adda <= "10101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101111";
				      t2adda <= "10101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110000";
				      t2adda <= "10110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000010111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110001";
				      t2adda <= "10110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110010";
				      t2adda <= "10110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110011";
				      t2adda <= "10110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110100";
				      t2adda <= "10110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000010111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110101";
				      t2adda <= "10110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000010111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110110";
				      t2adda <= "10110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110111";
				      t2adda <= "10110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111000";
				      t2adda <= "10111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111001";
				      t2adda <= "10111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111010";
				      t2adda <= "10111010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111011";
				      t2adda <= "10111011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111100";
				      t2adda <= "10111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111101";
				      t2adda <= "10111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111110";
				      t2adda <= "10111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111111";
				      t2adda <= "10111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000000";
				      t2adda <= "11000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000001";
				      t2adda <= "11000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000010";
				      t2adda <= "11000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000011";
				      t2adda <= "11000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000100";
				      t2adda <= "11000100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000101";
				      t2adda <= "11000101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000110";
				      t2adda <= "11000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000111";
				      t2adda <= "11000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001000";
				      t2adda <= "11001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001001";
				      t2adda <= "11001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001010";
				      t2adda <= "11001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001011";
				      t2adda <= "11001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001100";
				      t2adda <= "11001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001101";
				      t2adda <= "11001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001110";
				      t2adda <= "11001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001111";
				      t2adda <= "11001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010000";
				      t2adda <= "11010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010001";
				      t2adda <= "11010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010010";
				      t2adda <= "11010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010011";
				      t2adda <= "11010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010100";
				      t2adda <= "11010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010101";
				      t2adda <= "11010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010110";
				      t2adda <= "11010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010111";
				      t2adda <= "11010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011000";
				      t2adda <= "11011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011001";
				      t2adda <= "11011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011010";
				      t2adda <= "11011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011011";
				      t2adda <= "11011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011100";
				      t2adda <= "11011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011101";
				      t2adda <= "11011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011110";
				      t2adda <= "11011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011111";
				      t2adda <= "11011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100000";
				      t2adda <= "11100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100001";
				      t2adda <= "11100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100010";
				      t2adda <= "11100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100011";
				      t2adda <= "11100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100100";
				      t2adda <= "11100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100101";
				      t2adda <= "11100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100110";
				      t2adda <= "11100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100111";
				      t2adda <= "11100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101000";
				      t2adda <= "11101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101001";
				      t2adda <= "11101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101010";
				      t2adda <= "11101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101011";
				      t2adda <= "11101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101100";
				      t2adda <= "11101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101101";
				      t2adda <= "11101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101110";
				      t2adda <= "11101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101111";
				      t2adda <= "11101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110000";
				      t2adda <= "11110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000011111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110001";
				      t2adda <= "11110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110010";
				      t2adda <= "11110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110011";
				      t2adda <= "11110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110100";
				      t2adda <= "11110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000011111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110101";
				      t2adda <= "11110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000011111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110110";
				      t2adda <= "11110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110111";
				      t2adda <= "11110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111000";
				      t2adda <= "11111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000100000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111001";
				      t2adda <= "11111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="000100000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111010";
				      t2adda <= "11111010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="000100000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111011";
				      t2adda <= "11111011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="000100000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111100";
				      t2adda <= "11111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				                              
				elsif cntr1 ="000100000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111101";
				      t2adda <= "11111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000100000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111110";
				      t2adda <= "11111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                          
				                                          
				                                          
				elsif cntr1 ="000100001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111111";
				      t2adda <= "11111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                
				                                
				                                
				elsif cntr1 ="000100001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000000";
				      t2adda <= "00000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000100001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
				      t2adda <= "00000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
				      t2adda <= "00000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
				      t2adda <= "00000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000100";
				      t2adda <= "00000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
				      t2adda <= "00000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000111";
				      t2adda <= "00000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001000";
				      t2adda <= "00001000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000100010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001010";
				      t2adda <= "00001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
				      t2adda <= "00001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
				      t2adda <= "00001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
				      t2adda <= "00001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001111";
				      t2adda <= "00001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010000";
				      t2adda <= "00010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000100011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010001";
				      t2adda <= "00010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010010";
				      t2adda <= "00010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010011";
				      t2adda <= "00010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010100";
				      t2adda <= "00010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010101";
				      t2adda <= "00010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010110";
				      t2adda <= "00010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010111";
				      t2adda <= "00010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011000";
				      t2adda <= "00011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000100100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
				      t2adda <= "00011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011100";
				      t2adda <= "00011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011101";
				      t2adda <= "00011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011110";
				      t2adda <= "00011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011111";
				      t2adda <= "00011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100000";
				      t2adda <= "00100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000100101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100001";
				      t2adda <= "00100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
				      t2adda <= "00100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100110";
				      t2adda <= "00100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100111";
				      t2adda <= "00100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000100110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101001";
				      t2adda <= "00101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101010";
				      t2adda <= "00101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101011";
				      t2adda <= "00101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101100";
				      t2adda <= "00101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101101";
				      t2adda <= "00101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101110";
				      t2adda <= "00101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101111";
				      t2adda <= "00101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000100111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110000";
				      t2adda <= "00110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000100111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110001";
				      t2adda <= "00110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
				      t2adda <= "00110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
				      t2adda <= "00110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
				      t2adda <= "00110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
				      t2adda <= "00110110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111000";
				      t2adda <= "00111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
				      t2adda <= "00111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111010";
				      t2adda <= "00111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111011";
				      t2adda <= "00111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111100";
				      t2adda <= "00111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111101";
				      t2adda <= "00111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111110";
				      t2adda <= "00111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111111";
				      t2adda <= "00111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000000";
				      t2adda <= "01000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000101001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000001";
				      t2adda <= "01000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000010";
				      t2adda <= "01000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000011";
				      t2adda <= "01000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000100";
				      t2adda <= "01000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000101";
				      t2adda <= "01000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000110";
				      t2adda <= "01000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
				      t2adda <= "01000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001000";
				      t2adda <= "01001000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
				      t2adda <= "01001001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001010";
				      t2adda <= "01001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
				      t2adda <= "01001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001100";
				      t2adda <= "01001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001101";
				      t2adda <= "01001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001110";
				      t2adda <= "01001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001111";
				      t2adda <= "01001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010000";
				      t2adda <= "01010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000101011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010001";
				      t2adda <= "01010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
				      t2adda <= "01010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010011";
				      t2adda <= "01010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
				      t2adda <= "01010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
				      t2adda <= "01010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
				      t2adda <= "01010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
				      t2adda <= "01010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
				      t2adda <= "01011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011001";
				      t2adda <= "01011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
				      t2adda <= "01011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
				      t2adda <= "01011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
				      t2adda <= "01011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011101";
				      t2adda <= "01011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011110";
				      t2adda <= "01011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011111";
				      t2adda <= "01011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
				      t2adda <= "01100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000101101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100010";
				      t2adda <= "01100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100011";
				      t2adda <= "01100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100100";
				      t2adda <= "01100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100101";
				      t2adda <= "01100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100110";
				      t2adda <= "01100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100111";
				      t2adda <= "01100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
				      t2adda <= "01101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000101110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101001";
				      t2adda <= "01101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
				      t2adda <= "01101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
				      t2adda <= "01101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101101";
				      t2adda <= "01101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101110";
				      t2adda <= "01101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101111";
				      t2adda <= "01101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000101111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110000";
				      t2adda <= "01110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000101111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110001";
				      t2adda <= "01110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
				      t2adda <= "01110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110011";
				      t2adda <= "01110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110100";
				      t2adda <= "01110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110101";
				      t2adda <= "01110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110110";
				      t2adda <= "01110110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110111";
				      t2adda <= "01110111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111000";
				      t2adda <= "01111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111001";
				      t2adda <= "01111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="000110000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111010";
				      t2adda <= "01111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				elsif cntr1 ="000110000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111011";
				      t2adda <= "01111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				elsif cntr1 ="000110000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111100";
				      t2adda <= "01111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				                              
				elsif cntr1 ="000110000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111101";
				      t2adda <= "01111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000110000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111110";
				      t2adda <= "01111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                        
				                                        
				                                        
				elsif cntr1 ="000110001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111111";
				      t2adda <= "01111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                      
				                                      
				                                      
				elsif cntr1 ="000110001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000000";
				      t2adda <= "10000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000001";
				      t2adda <= "10000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000010";
				      t2adda <= "10000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000011";
				      t2adda <= "10000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000100";
				      t2adda <= "10000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000101";
				      t2adda <= "10000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000110";
				      t2adda <= "10000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000111";
				      t2adda <= "10000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001000";
				      t2adda <= "10001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000110010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001001";
				      t2adda <= "10001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001010";
				      t2adda <= "10001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001011";
				      t2adda <= "10001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001100";
				      t2adda <= "10001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001101";
				      t2adda <= "10001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001110";
				      t2adda <= "10001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001111";
				      t2adda <= "10001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010000";
				      t2adda <= "10010000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010001";
				      t2adda <= "10010001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010010";
				      t2adda <= "10010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010011";
				      t2adda <= "10010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010100";
				      t2adda <= "10010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010101";
				      t2adda <= "10010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010110";
				      t2adda <= "10010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010111";
				      t2adda <= "10010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011000";
				      t2adda <= "10011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000110100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011001";
				      t2adda <= "10011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011010";
				      t2adda <= "10011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011011";
				      t2adda <= "10011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011100";
				      t2adda <= "10011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011101";
				      t2adda <= "10011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011110";
				      t2adda <= "10011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011111";
				      t2adda <= "10011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100000";
				      t2adda <= "10100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100001";
				      t2adda <= "10100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100010";
				      t2adda <= "10100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100011";
				      t2adda <= "10100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100100";
				      t2adda <= "10100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100101";
				      t2adda <= "10100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100110";
				      t2adda <= "10100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100111";
				      t2adda <= "10100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101000";
				      t2adda <= "10101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000110110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101001";
				      t2adda <= "10101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101010";
				      t2adda <= "10101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101011";
				      t2adda <= "10101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101100";
				      t2adda <= "10101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101101";
				      t2adda <= "10101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101110";
				      t2adda <= "10101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101111";
				      t2adda <= "10101111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110000";
				      t2adda <= "10110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110001";
				      t2adda <= "10110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110010";
				      t2adda <= "10110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110011";
				      t2adda <= "10110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110100";
				      t2adda <= "10110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110101";
				      t2adda <= "10110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000110111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110110";
				      t2adda <= "10110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110111";
				      t2adda <= "10110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111000";
				      t2adda <= "10111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111001";
				      t2adda <= "10111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111010";
				      t2adda <= "10111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111011";
				      t2adda <= "10111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111100";
				      t2adda <= "10111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111101";
				      t2adda <= "10111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111110";
				      t2adda <= "10111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111111";
				      t2adda <= "10111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000000";
				      t2adda <= "11000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000001";
				      t2adda <= "11000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000010";
				      t2adda <= "11000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000011";
				      t2adda <= "11000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000100";
				      t2adda <= "11000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000101";
				      t2adda <= "11000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000110";
				      t2adda <= "11000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000111";
				      t2adda <= "11000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001000";
				      t2adda <= "11001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000111010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001001";
				      t2adda <= "11001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001010";
				      t2adda <= "11001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001011";
				      t2adda <= "11001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001100";
				      t2adda <= "11001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001101";
				      t2adda <= "11001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001110";
				      t2adda <= "11001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001111";
				      t2adda <= "11001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010000";
				      t2adda <= "11010000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010001";
				      t2adda <= "11010001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010010";
				      t2adda <= "11010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010011";
				      t2adda <= "11010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010100";
				      t2adda <= "11010100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010101";
				      t2adda <= "11010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010110";
				      t2adda <= "11010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010111";
				      t2adda <= "11010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011000";
				      t2adda <= "11011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="000111100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011001";
				      t2adda <= "11011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011010";
				      t2adda <= "11011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011011";
				      t2adda <= "11011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011100";
				      t2adda <= "11011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011101";
				      t2adda <= "11011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011110";
				      t2adda <= "11011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011111";
				      t2adda <= "11011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100000";
				      t2adda <= "11100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100001";
				      t2adda <= "11100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100010";
				      t2adda <= "11100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100011";
				      t2adda <= "11100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100100";
				      t2adda <= "11100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100101";
				      t2adda <= "11100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100110";
				      t2adda <= "11100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100111";
				      t2adda <= "11100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101000";
				      t2adda <= "11101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="000111110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101001";
				      t2adda <= "11101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101010";
				      t2adda <= "11101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101011";
				      t2adda <= "11101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101100";
				      t2adda <= "11101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101101";
				      t2adda <= "11101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101110";
				      t2adda <= "11101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101111";
				      t2adda <= "11101111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110000";
				      t2adda <= "11110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110001";
				      t2adda <= "11110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110010";
				      t2adda <= "11110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110011";
				      t2adda <= "11110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110100";
				      t2adda <= "11110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110101";
				      t2adda <= "11110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="000111111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110110";
				      t2adda <= "11110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110111";
				      t2adda <= "11110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111000";
				      t2adda <= "11111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="001000000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111001";
				      t2adda <= "11111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="001000000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111010";
				      t2adda <= "11111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				elsif cntr1 ="001000000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111011";
				      t2adda <= "11111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				elsif cntr1 ="001000000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111100";
				      t2adda <= "11111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				                              
				elsif cntr1 ="001000000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111101";
				      t2adda <= "11111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001000000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111110";
				      t2adda <= "11111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                         
				                                         
				                                         
				elsif cntr1 ="001000001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111111";
				      t2adda <= "11111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                  
				                                  
				                                  
				elsif cntr1 ="001000001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000000";
				      t2adda <= "00000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000001";
				      t2adda <= "00000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000010";
				      t2adda <= "00000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000011";
				      t2adda <= "00000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000100";
				      t2adda <= "00000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000101";
				      t2adda <= "00000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000110";
				      t2adda <= "00000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00000111";
				      t2adda <= "00000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001000";
				      t2adda <= "00001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001001";
				      t2adda <= "00001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001010";
				      t2adda <= "00001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001011";
				      t2adda <= "00001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001100";
				      t2adda <= "00001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001101";
				      t2adda <= "00001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001110";
				      t2adda <= "00001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00001111";
				      t2adda <= "00001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010000";
				      t2adda <= "00010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010001";
				      t2adda <= "00010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010010";
				      t2adda <= "00010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010011";
				      t2adda <= "00010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010100";
				      t2adda <= "00010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010101";
				      t2adda <= "00010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010110";
				      t2adda <= "00010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00010111";
				      t2adda <= "00010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011000";
				      t2adda <= "00011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001000100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011001";
				      t2adda <= "00011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011010";
				      t2adda <= "00011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011011";
				      t2adda <= "00011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011100";
				      t2adda <= "00011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011101";
				      t2adda <= "00011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011110";
				      t2adda <= "00011110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00011111";
				      t2adda <= "00011111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100000";
				      t2adda <= "00100000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100001";
				      t2adda <= "00100001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100010";
				      t2adda <= "00100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100011";
				      t2adda <= "00100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100100";
				      t2adda <= "00100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100101";
				      t2adda <= "00100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100110";
				      t2adda <= "00100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00100111";
				      t2adda <= "00100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101000";
				      t2adda <= "00101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101001";
				      t2adda <= "00101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101010";
				      t2adda <= "00101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101011";
				      t2adda <= "00101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101100";
				      t2adda <= "00101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101101";
				      t2adda <= "00101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101110";
				      t2adda <= "00101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00101111";
				      t2adda <= "00101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110000";
				      t2adda <= "00110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110001";
				      t2adda <= "00110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110010";
				      t2adda <= "00110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110011";
				      t2adda <= "00110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110100";
				      t2adda <= "00110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110101";
				      t2adda <= "00110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001000111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110110";
				      t2adda <= "00110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00110111";
				      t2adda <= "00110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111000";
				      t2adda <= "00111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="001001000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111001";
				      t2adda <= "00111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111010";
				      t2adda <= "00111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111011";
				      t2adda <= "00111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111100";
				      t2adda <= "00111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111101";
				      t2adda <= "00111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111110";
				      t2adda <= "00111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "00111111";
				      t2adda <= "00111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001001001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000000";
				      t2adda <= "01000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000001";
				      t2adda <= "01000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000010";
				      t2adda <= "01000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000011";
				      t2adda <= "01000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000100";
				      t2adda <= "01000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000101";
				      t2adda <= "01000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000110";
				      t2adda <= "01000110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01000111";
				      t2adda <= "01000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001000";
				      t2adda <= "01001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001001";
				      t2adda <= "01001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001010";
				      t2adda <= "01001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001011";
				      t2adda <= "01001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001100";
				      t2adda <= "01001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001101";
				      t2adda <= "01001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001110";
				      t2adda <= "01001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01001111";
				      t2adda <= "01001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010000";
				      t2adda <= "01010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010001";
				      t2adda <= "01010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010010";
				      t2adda <= "01010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010011";
				      t2adda <= "01010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010100";
				      t2adda <= "01010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010101";
				      t2adda <= "01010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010110";
				      t2adda <= "01010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01010111";
				      t2adda <= "01010111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011000";
				      t2adda <= "01011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001001100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011001";
				      t2adda <= "01011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011010";
				      t2adda <= "01011010";
						t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011011";
				      t2adda <= "01011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011100";
				      t2adda <= "01011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011101";
				      t2adda <= "01011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011110";
				      t2adda <= "01011110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01011111";
				      t2adda <= "01011111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100000";
				      t2adda <= "01100000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101010" THEN
				      
				      
						t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100001";
				      t2adda <= "01100001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100010";
				      t2adda <= "01100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100011";
				      t2adda <= "01100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100100";
				      t2adda <= "01100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
						
				      
				elsif cntr1 ="001001101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100101";
				      t2adda <= "01100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100110";
				      t2adda <= "01100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01100111";
				      t2adda <= "01100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101000";
				      t2adda <= "01101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101001";
				      t2adda <= "01101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101010";
				      t2adda <= "01101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101011";
						t2adda <= "01101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101100";
				      t2adda <= "01101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101101";
				      t2adda <= "01101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101110";
				      t2adda <= "01101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01101111";
				      t2adda <= "01101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110000";
				      t2adda <= "01110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110001";
				      t2adda <= "01110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111011" THEN
				      
						
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110010";
				      t2adda <= "01110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110011";
				      t2adda <= "01110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110100";
				      t2adda <= "01110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001001111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110101";
				      t2adda <= "01110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
						
				      
				      
				elsif cntr1 ="001001111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110110";
				      t2adda <= "01110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01110111";
				      t2adda <= "01110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111000";
				      t2adda <= "01111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="001010000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111001";
				      t2adda <= "01111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="001010000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111010";
				      t2adda <= "01111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				elsif cntr1 ="001010000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111011";
				      t2adda <= "01111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				elsif cntr1 ="001010000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
					  t1adda <= "01111100";
				      t2adda <= "01111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				                              
				elsif cntr1 ="001010000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111101";
				      t2adda <= "01111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001010000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111110";
				      t2adda <= "01111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                       
				                                       
				                                       
				elsif cntr1 ="001010001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "01111111";
				      t2adda <= "01111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                         
				                                         
				                                         
				elsif cntr1 ="001010001001" THEN
				
				
					  t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000000";
				      t2adda <= "10000000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000001";
				      t2adda <= "10000001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000010";
				      t2adda <= "10000010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001100" THEN
						
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000011";
				      t2adda <= "10000011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000100";
				      t2adda <= "10000100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000101";
				      t2adda <= "10000101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000110";
				      t2adda <= "10000110";
				      t1dina <= bfrjout;
						t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10000111";
				      t2adda <= "10000111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001000";
				      t2adda <= "10001000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001001";
				      t2adda <= "10001001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001010";
				      t2adda <= "10001010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001011";
				      t2adda <= "10001011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001100";
				      t2adda <= "10001100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010110" THEN
				      
				      
				      t1wea <= '1';
						t2wea <= '1';
				      t1adda <= "10001101";
				      t2adda <= "10001101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001110";
				      t2adda <= "10001110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10001111";
				      t2adda <= "10001111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010000";
				      t2adda <= "10010000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
						
				elsif cntr1 ="001010011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010001";
				      t2adda <= "10010001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010010";
				      t2adda <= "10010010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010011";
				      t2adda <= "10010011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010100";
				      t2adda <= "10010100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010101";
				      t2adda <= "10010101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010110";
				      t2adda <= "10010110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10010111";
				      t2adda <= "10010111";
						t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011000";
				      t2adda <= "10011000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011001";
				      t2adda <= "10011001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011010";
				      t2adda <= "10011010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011011";
				      t2adda <= "10011011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011100";
				      t2adda <= "10011100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011101";
				      t2adda <= "10011101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010100111" THEN
				      
				      
						t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011110";
				      t2adda <= "10011110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10011111";
				      t2adda <= "10011111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100000";
				      t2adda <= "10100000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100001";
				      t2adda <= "10100001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
						
				      
				elsif cntr1 ="001010101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100010";
				      t2adda <= "10100010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100011";
				      t2adda <= "10100011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100100";
				      t2adda <= "10100100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100101";
				      t2adda <= "10100101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100110";
				      t2adda <= "10100110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10100111";
				      t2adda <= "10100111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101000";
						t2adda <= "10101000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101001";
				      t2adda <= "10101001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101010";
				      t2adda <= "10101010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101011";
				      t2adda <= "10101011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101100";
				      t2adda <= "10101100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101101";
				      t2adda <= "10101101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101110";
				      t2adda <= "10101110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111000" THEN
				      
						
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10101111";
				      t2adda <= "10101111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110000";
				      t2adda <= "10110000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110001";
				      t2adda <= "10110001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110010";
				      t2adda <= "10110010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
						
				      
				      
				elsif cntr1 ="001010111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110011";
				      t2adda <= "10110011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110100";
				      t2adda <= "10110100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110101";
				      t2adda <= "10110101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110110";
				      t2adda <= "10110110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10110111";
				      t2adda <= "10110111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111000";
				      t2adda <= "10111000";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				elsif cntr1 ="001011000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
						t1adda <= "10111001";
				      t2adda <= "10111001";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111010";
				      t2adda <= "10111010";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111011";
				      t2adda <= "10111011";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111100";
				      t2adda <= "10111100";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111101";
				      t2adda <= "10111101";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111110";
				      t2adda <= "10111110";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "10111111";
				      t2adda <= "10111111";
				      t1dina <= bfrjout;
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001011001001" THEN
						
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000000";
				      t2adda <= "11000000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000001";
				      t2adda <= "11000001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000010";
				      t2adda <= "11000010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000011";
				      t2adda <= "11000011";
				      t1dina <= bfrjplout;
						t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000100";
				      t2adda <= "11000100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000101";
				      t2adda <= "11000101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000110";
				      t2adda <= "11000110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11000111";
				      t2adda <= "11000111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001000";
				      t2adda <= "11001000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001001";
				      t2adda <= "11001001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010011" THEN
				      
				      
				      t1wea <= '1';
						t2wea <= '1';
				      t1adda <= "11001010";
				      t2adda <= "11001010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001011";
				      t2adda <= "11001011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001100";
				      t2adda <= "11001100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001101";
				      t2adda <= "11001101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
						
				elsif cntr1 ="001011010111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001110";
				      t2adda <= "11001110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11001111";
				      t2adda <= "11001111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010000";
				      t2adda <= "11010000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010001";
				      t2adda <= "11010001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010010";
				      t2adda <= "11010010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010011";
				      t2adda <= "11010011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010100";
				      t2adda <= "11010100";
						t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010101";
				      t2adda <= "11010101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010110";
				      t2adda <= "11010110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11010111";
				      t2adda <= "11010111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011000";
				      t2adda <= "11011000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011001";
				      t2adda <= "11011001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011010";
				      t2adda <= "11011010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100100" THEN
				      
				      
						t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011011";
				      t2adda <= "11011011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011100";
				      t2adda <= "11011100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011101";
				      t2adda <= "11011101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011110";
				      t2adda <= "11011110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
						
				      
				elsif cntr1 ="001011101000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11011111";
				      t2adda <= "11011111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100000";
				      t2adda <= "11100000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100001";
				      t2adda <= "11100001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100010";
				      t2adda <= "11100010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100011";
				      t2adda <= "11100011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100100";
				      t2adda <= "11100100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100101";
						t2adda <= "11100101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100110";
				      t2adda <= "11100110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11100111";
				      t2adda <= "11100111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101000";
				      t2adda <= "11101000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101001";
				      t2adda <= "11101001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101010";
				      t2adda <= "11101010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101011";
				      t2adda <= "11101011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110101" THEN
				      
						
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101100";
				      t2adda <= "11101100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101101";
				      t2adda <= "11101101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101110";
				      t2adda <= "11101110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11101111";
				      t2adda <= "11101111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
						
				      
				      
				elsif cntr1 ="001011111001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110000";
				      t2adda <= "11110000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110001";
				      t2adda <= "11110001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110010";
				      t2adda <= "11110010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110011";
				      t2adda <= "11110011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110100";
				      t2adda <= "11110100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111110" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11110101";
				      t2adda <= "11110101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
						t1adda <= "11110110";
				      t2adda <= "11110110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
						t1adda <= "11110111";
				      t2adda <= "11110111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000001" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
						t1adda <= "11111000";
				      t2adda <= "11111000";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				      
				      
				elsif cntr1 ="001100000010" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111001";
				      t2adda <= "11111001";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				            
				            
				            
				elsif cntr1 ="001100000011" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111010";
				      t2adda <= "11111010";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                  
				                  
				                  
				elsif cntr1 ="001100000100" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111011";
				      t2adda <= "11111011";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                        
				                        
				                        
				elsif cntr1 ="001100000101" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111100";
				      t2adda <= "11111100";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                              
				                              
				                              
				elsif cntr1 ="001100000110" THEN
						
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111101";
				      t2adda <= "11111101";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                    
				                                    
				                                    
				 elsif cntr1 ="001100000111" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111110";
				      t2adda <= "11111110";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                          
				                                          
				                                          
				 elsif cntr1 ="001100001000" THEN
				      
				      
				      t1wea <= '1';
				      t2wea <= '1';
				      t1adda <= "11111111";
				      t2adda <= "11111111";
				      t1dina <= bfrjplout;
				      t2dina <= bfrjout;
				                                          
				                                          
				                                          
				elsif cntr1 ="001100001001" THEN
				
				
					  t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000000";
				      ioaddb <= "010000000";
				      t1dina <= bfrjout;
						iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000001";
				      ioaddb <= "010000001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000010";
				      ioaddb <= "010000010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000011";
				      ioaddb <= "010000011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000100";
				      ioaddb <= "010000100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000101";
				      ioaddb <= "010000101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100001111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00000110";
				      ioaddb <= "010000110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010000" THEN
				      
				      
				      t1wea <= '1';
						ioweb <= '1';
				      t1adda <= "00000111";
				      ioaddb <= "010000111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001000";
				      ioaddb <= "010001000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001001";
				      ioaddb <= "010001001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001010";
				      ioaddb <= "010001010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
						
				elsif cntr1 ="001100010100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001011";
				      ioaddb <= "010001011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001100";
				      ioaddb <= "010001100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001101";
				      ioaddb <= "010001101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100010111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001110";
				      ioaddb <= "010001110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00001111";
				      ioaddb <= "010001111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010000";
				      ioaddb <= "010010000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010001";
				      ioaddb <= "010010001";
						t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010010";
				      ioaddb <= "010010010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010011";
				      ioaddb <= "010010011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010100";
				      ioaddb <= "010010100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010101";
				      ioaddb <= "010010101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100011111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010110";
				      ioaddb <= "010010110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00010111";
				      ioaddb <= "010010111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100001" THEN
				      
				      
						t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011000";
				      ioaddb <= "010011000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011001";
				      ioaddb <= "010011001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011010";
				      ioaddb <= "010011010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011011";
				      ioaddb <= "010011011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
						
				      
				elsif cntr1 ="001100100101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011100";
				      ioaddb <= "010011100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011101";
				      ioaddb <= "010011101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100100111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011110";
				      ioaddb <= "010011110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00011111";
				      ioaddb <= "010011111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100000";
				      ioaddb <= "010100000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100001";
				      ioaddb <= "010100001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100010";
						ioaddb <= "010100010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100011";
				      ioaddb <= "010100011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100100";
				      ioaddb <= "010100100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100101";
				      ioaddb <= "010100101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100101111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100110";
				      ioaddb <= "010100110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00100111";
				      ioaddb <= "010100111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101000";
				      ioaddb <= "010101000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110010" THEN
				      
						
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101001";
				      ioaddb <= "010101001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101010";
				      ioaddb <= "010101010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101011";
				      ioaddb <= "010101011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101100";
				      ioaddb <= "010101100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
						
				      
				      
				elsif cntr1 ="001100110110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101101";
				      ioaddb <= "010101101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100110111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101110";
				      ioaddb <= "010101110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00101111";
				      ioaddb <= "010101111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110000";
				      ioaddb <= "010110000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110001";
				      ioaddb <= "010110001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110010";
				      ioaddb <= "010110010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
						t1adda <= "00110011";
				      ioaddb <= "010110011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110100";
				      ioaddb <= "010110100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110101";
				      ioaddb <= "010110101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001100111111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110110";
				      ioaddb <= "010110110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00110111";
				      ioaddb <= "010110111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111000";
				      ioaddb <= "010111000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111001";
				      ioaddb <= "010111001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000011" THEN
						
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111010";
				      ioaddb <= "010111010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111011";
				      ioaddb <= "010111011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111100";
				      ioaddb <= "010111100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111101";
				      ioaddb <= "010111101";
				      t1dina <= bfrjout;
						iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101000111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111110";
				      ioaddb <= "010111110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "00111111";
				      ioaddb <= "010111111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000000";
				      ioaddb <= "011000000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000001";
				      ioaddb <= "011000001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000010";
				      ioaddb <= "011000010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000011";
				      ioaddb <= "011000011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001101" THEN
				      
				      
				      t1wea <= '1';
						ioweb <= '1';
				      t1adda <= "01000100";
				      ioaddb <= "011000100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000101";
				      ioaddb <= "011000101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101001111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000110";
				      ioaddb <= "011000110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01000111";
				      ioaddb <= "011000111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
						
				elsif cntr1 ="001101010001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001000";
				      ioaddb <= "011001000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001001";
				      ioaddb <= "011001001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001010";
				      ioaddb <= "011001010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001011";
				      ioaddb <= "011001011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001100";
				      ioaddb <= "011001100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001101";
				      ioaddb <= "011001101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101010111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001110";
				      ioaddb <= "011001110";
						t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01001111";
				      ioaddb <= "011001111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010000";
				      ioaddb <= "011010000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010001";
				      ioaddb <= "011010001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010010";
				      ioaddb <= "011010010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010011";
				      ioaddb <= "011010011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010100";
				      ioaddb <= "011010100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011110" THEN
				      
				      
						t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010101";
				      ioaddb <= "011010101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101011111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010110";
				      ioaddb <= "011010110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01010111";
				      ioaddb <= "011010111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011000";
				      ioaddb <= "011011000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
						
				      
				elsif cntr1 ="001101100010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011001";
				      ioaddb <= "011011001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011010";
				      ioaddb <= "011011010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011011";
				      ioaddb <= "011011011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011100";
				      ioaddb <= "011011100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011101";
				      ioaddb <= "011011101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101100111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011110";
				      ioaddb <= "011011110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01011111";
						ioaddb <= "011011111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100000";
				      ioaddb <= "011100000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100001";
				      ioaddb <= "011100001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100010";
				      ioaddb <= "011100010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100011";
				      ioaddb <= "011100011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100100";
				      ioaddb <= "011100100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100101";
				      ioaddb <= "011100101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101101111" THEN
				      
						
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100110";
				      ioaddb <= "011100110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01100111";
				      ioaddb <= "011100111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101000";
				      ioaddb <= "011101000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101001";
				      ioaddb <= "011101001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
						
				      
				      
				elsif cntr1 ="001101110011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101010";
				      ioaddb <= "011101010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101011";
				      ioaddb <= "011101011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101100";
				      ioaddb <= "011101100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101101";
				      ioaddb <= "011101101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101110111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101110";
				      ioaddb <= "011101110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01101111";
				      ioaddb <= "011101111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111001" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
						t1adda <= "01110000";
				      ioaddb <= "011110000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110001";
				      ioaddb <= "011110001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110010";
				      ioaddb <= "011110010";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110011";
				      ioaddb <= "011110011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110100";
				      ioaddb <= "011110100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110101";
				      ioaddb <= "011110101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001101111111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110110";
				      ioaddb <= "011110110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110000000" THEN
						
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01110111";
				      ioaddb <= "011110111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110000001" THEN
						
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111000";
				      ioaddb <= "011111000";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				      
				      
				elsif cntr1 ="001110000010" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111001";
				      ioaddb <= "011111001";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="001110000011" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111010";
				      ioaddb <= "011111010";
				      t1dina <= bfrjout;
						iodinb <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="001110000100" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111011";
				      ioaddb <= "011111011";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="001110000101" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111100";
				      ioaddb <= "011111100";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="001110000110" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111101";
				      ioaddb <= "011111101";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001110000111" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111110";
				      ioaddb <= "011111110";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				                                          
				                                          
				                                          
				elsif cntr1 ="001110001000" THEN
				      
				      
				      t1wea <= '1';
				      ioweb <= '1';
				      t1adda <= "01111111";
				      ioaddb <= "011111111";
				      t1dina <= bfrjout;
				      iodinb <= bfrjplout;
				                                   
				                                   
				                                   
				elsif cntr1 ="001110001001" THEN
				
				
					  
				      ioweb <= '1';
				      
				      ioaddb <= "000000000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110001010" THEN
				      
				      
				      
					  ioweb <= '1';
				      
				      ioaddb <= "000000001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000100";
				      
				      iodinb <= bfrjplout;
				      
				      
						
				elsif cntr1 ="001110001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001011";
						
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011011" THEN
				      
				      
						
				      ioweb <= '1';
				      
				      ioaddb <= "000010010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010101";
				      
				      iodinb <= bfrjplout;
				      
						
				      
				elsif cntr1 ="001110011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
						ioaddb <= "000011100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101100" THEN
				      
						
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100110";
				      
				      iodinb <= bfrjplout;
						
				      
				      
				elsif cntr1 ="001110110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110110" THEN
				      
				      
				      
				      ioweb <= '1';
						
				      ioaddb <= "000101101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111101" THEN
						
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001110111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110111";
				      
						iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111000111" THEN
				      
				      
				      
						ioweb <= '1';
				      
				      ioaddb <= "000111110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000001";
				      
				      iodinb <= bfrjplout;
				      
				      
						
				elsif cntr1 ="001111001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001000";
						
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011000" THEN
				      
				      
						
				      ioweb <= '1';
				      
				      ioaddb <= "001001111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010010";
				      
				      iodinb <= bfrjplout;
				      
						
				      
				elsif cntr1 ="001111011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
						ioaddb <= "001011001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101001" THEN
				      
						
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100011";
				      
				      iodinb <= bfrjplout;
						
				      
				      
				elsif cntr1 ="001111101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110011" THEN
				      
				      
				      
				      ioweb <= '1';
						
				      ioaddb <= "001101010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101100";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111010" THEN
						
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110001";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110010";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110011";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110100";
				      
						iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110101";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001111111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110110";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="010000000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110111";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="010000000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111000";
				      
				      iodinb <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="010000000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111001";
				      
				      iodinb <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="010000000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111010";
				      
				      iodinb <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="010000000100" THEN
				      
				      
				      
						ioweb <= '1';
				      
				      ioaddb <= "001111011";
				      
				      iodinb <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="010000000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111100";
				      
				      iodinb <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="010000000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111101";
				      
				      iodinb <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="010000000111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111110";
				      
				      iodinb <= bfrjplout;
				                                        
				                                        
				                                  		
				elsif cntr1 ="010000001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111111";
				      
				      iodinb <= bfrjplout;
				                                    
				       
					
				                                  	
				elsif cntr1 ="010000001001" THEN
				
				elsif cntr1 ="010000001010" THEN
				
				
				
				
				
				
				
				
				
	
				
				END IF;					
			
			
			
			
			
			
			
			
			
			
			
				
				
			
				
				
			
			ELSIF cur_st = topwm THEN
			





				if cntr ="000000000000" THEN	
				      ioadda <= "000000001";
				      ioaddb <= "100000001";
				      
				      bfmod <= "01";
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000001";
				elsif cntr ="000000000001" THEN
				      ioadda <= "000000011";
				      ioaddb <= "100000011";
				      
				      
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000010";
				elsif cntr ="000000000010" THEN
				      ioadda <= "000000101";
				      ioaddb <= "100000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000011";
				elsif cntr ="000000000011" THEN
				      ioadda <= "000000111";
				      ioaddb <= "100000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000100";
				elsif cntr ="000000000100" THEN
				      ioadda <= "000001001";
				      ioaddb <= "100001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000101";
				elsif cntr ="000000000101" THEN
				      ioadda <= "000001011";
				      ioaddb <= "100001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000110";
				elsif cntr ="000000000110" THEN
				      ioadda <= "000001101";
				      ioaddb <= "100001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000000111";
				elsif cntr ="000000000111" THEN
				      ioadda <= "000001111";
				      ioaddb <= "100001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "000000001000";
				elsif cntr ="000000001000" THEN
				      ioadda <= "000010001";
				      ioaddb <= "100010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				      
				      
				      
				      cntr <= "000000001001";
				elsif cntr ="000000001001" THEN
				      ioadda <= "000010011";
				      ioaddb <= "100010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001010";
				elsif cntr ="000000001010" THEN
				      ioadda <= "000010101";
				      ioaddb <= "100010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001011";
				elsif cntr ="000000001011" THEN
				      ioadda <= "000010111";
				      ioaddb <= "100010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001100";
				elsif cntr ="000000001100" THEN
				      ioadda <= "000011001";
				      ioaddb <= "100011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001101";
				elsif cntr ="000000001101" THEN
				      ioadda <= "000011011";
				      ioaddb <= "100011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001110";
				elsif cntr ="000000001110" THEN
				      ioadda <= "000011101";
				      ioaddb <= "100011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000001111";
				elsif cntr ="000000001111" THEN
				      ioadda <= "000011111";
				      ioaddb <= "100011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010000";
				elsif cntr ="000000010000" THEN
				      ioadda <= "000100001";
				      ioaddb <= "100100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010001";
				elsif cntr ="000000010001" THEN
				      ioadda <= "000100011";
				      ioaddb <= "100100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010010";
				elsif cntr ="000000010010" THEN
				      ioadda <= "000100101";
				      ioaddb <= "100100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010011";
				elsif cntr ="000000010011" THEN
				      ioadda <= "000100111";
				      ioaddb <= "100100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010100";
				elsif cntr ="000000010100" THEN
				      ioadda <= "000101001";
				      ioaddb <= "100101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010101";
				elsif cntr ="000000010101" THEN
				      ioadda <= "000101011";
				      ioaddb <= "100101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010110";
				elsif cntr ="000000010110" THEN
				      ioadda <= "000101101";
				      ioaddb <= "100101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000010111";
				elsif cntr ="000000010111" THEN
				      ioadda <= "000101111";
				      ioaddb <= "100101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011000";
				elsif cntr ="000000011000" THEN
				      ioadda <= "000110001";
				      ioaddb <= "100110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011001";
				elsif cntr ="000000011001" THEN
				      ioadda <= "000110011";
				      ioaddb <= "100110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011010";
				elsif cntr ="000000011010" THEN
				      ioadda <= "000110101";
				      ioaddb <= "100110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011011";
				elsif cntr ="000000011011" THEN
				      ioadda <= "000110111";
				      ioaddb <= "100110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011100";
				elsif cntr ="000000011100" THEN
				      ioadda <= "000111001";
				      ioaddb <= "100111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011101";
				elsif cntr ="000000011101" THEN
				      ioadda <= "000111011";
				      ioaddb <= "100111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011110";
				elsif cntr ="000000011110" THEN
				      ioadda <= "000111101";
				      ioaddb <= "100111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000011111";
				elsif cntr ="000000011111" THEN
				      ioadda <= "000111111";
				      ioaddb <= "100111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100000";
				elsif cntr ="000000100000" THEN
				      ioadda <= "001000001";
				      ioaddb <= "101000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100001";
				elsif cntr ="000000100001" THEN
				      ioadda <= "001000011";
				      ioaddb <= "101000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100010";
				elsif cntr ="000000100010" THEN
				      ioadda <= "001000101";
				      ioaddb <= "101000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100011";
				elsif cntr ="000000100011" THEN
				      ioadda <= "001000111";
				      ioaddb <= "101000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100100";
				elsif cntr ="000000100100" THEN
				      ioadda <= "001001001";
				      ioaddb <= "101001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100101";
				elsif cntr ="000000100101" THEN
				      ioadda <= "001001011";
				      ioaddb <= "101001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100110";
				elsif cntr ="000000100110" THEN
				      ioadda <= "001001101";
				      ioaddb <= "101001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000100111";
				elsif cntr ="000000100111" THEN
				      ioadda <= "001001111";
				      ioaddb <= "101001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101000";
				elsif cntr ="000000101000" THEN
				      ioadda <= "001010001";
				      ioaddb <= "101010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101001";
				elsif cntr ="000000101001" THEN
				      ioadda <= "001010011";
				      ioaddb <= "101010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101010";
				elsif cntr ="000000101010" THEN
				      ioadda <= "001010101";
				      ioaddb <= "101010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101011";
				elsif cntr ="000000101011" THEN
				      ioadda <= "001010111";
				      ioaddb <= "101010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101100";
				elsif cntr ="000000101100" THEN
				      ioadda <= "001011001";
				      ioaddb <= "101011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101101";
				elsif cntr ="000000101101" THEN
				      ioadda <= "001011011";
				      ioaddb <= "101011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101110";
				elsif cntr ="000000101110" THEN
				      ioadda <= "001011101";
				      ioaddb <= "101011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000101111";
				elsif cntr ="000000101111" THEN
				      ioadda <= "001011111";
				      ioaddb <= "101011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110000";
				elsif cntr ="000000110000" THEN
				      ioadda <= "001100001";
				      ioaddb <= "101100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110001";
				elsif cntr ="000000110001" THEN
				      ioadda <= "001100011";
				      ioaddb <= "101100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110010";
				elsif cntr ="000000110010" THEN
				      ioadda <= "001100101";
				      ioaddb <= "101100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110011";
				elsif cntr ="000000110011" THEN
				      ioadda <= "001100111";
				      ioaddb <= "101100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110100";
				elsif cntr ="000000110100" THEN
				      ioadda <= "001101001";
				      ioaddb <= "101101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110101";
				elsif cntr ="000000110101" THEN
				      ioadda <= "001101011";
				      ioaddb <= "101101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110110";
				elsif cntr ="000000110110" THEN
				      ioadda <= "001101101";
				      ioaddb <= "101101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000110111";
				elsif cntr ="000000110111" THEN
				      ioadda <= "001101111";
				      ioaddb <= "101101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111000";
				elsif cntr ="000000111000" THEN
				      ioadda <= "001110001";
				      ioaddb <= "101110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111001";
				elsif cntr ="000000111001" THEN
				      ioadda <= "001110011";
				      ioaddb <= "101110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111010";
				elsif cntr ="000000111010" THEN
				      ioadda <= "001110101";
				      ioaddb <= "101110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111011";
				elsif cntr ="000000111011" THEN
				      ioadda <= "001110111";
				      ioaddb <= "101110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111100";
				elsif cntr ="000000111100" THEN
				      ioadda <= "001111001";
				      ioaddb <= "101111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111101";
				elsif cntr ="000000111101" THEN
				      ioadda <= "001111011";
				      ioaddb <= "101111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111110";
				elsif cntr ="000000111110" THEN
				      ioadda <= "001111101";
				      ioaddb <= "101111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000000111111";
				elsif cntr ="000000111111" THEN
				      ioadda <= "001111111";
				      ioaddb <= "101111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000000";
				elsif cntr ="000001000000" THEN
				      ioadda <= "010000001";
				      ioaddb <= "110000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000001";
				elsif cntr ="000001000001" THEN
				      ioadda <= "010000011";
				      ioaddb <= "110000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000010";
				elsif cntr ="000001000010" THEN
				      ioadda <= "010000101";
				      ioaddb <= "110000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000011";
				elsif cntr ="000001000011" THEN
				      ioadda <= "010000111";
				      ioaddb <= "110000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000100";
				elsif cntr ="000001000100" THEN
				      ioadda <= "010001001";
				      ioaddb <= "110001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000101";
				elsif cntr ="000001000101" THEN
				      ioadda <= "010001011";
				      ioaddb <= "110001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000110";
				elsif cntr ="000001000110" THEN
				      ioadda <= "010001101";
				      ioaddb <= "110001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001000111";
				elsif cntr ="000001000111" THEN
				      ioadda <= "010001111";
				      ioaddb <= "110001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001000";
				elsif cntr ="000001001000" THEN
				      ioadda <= "010010001";
				      ioaddb <= "110010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001001";
				elsif cntr ="000001001001" THEN
				      ioadda <= "010010011";
				      ioaddb <= "110010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001010";
				elsif cntr ="000001001010" THEN
				      ioadda <= "010010101";
				      ioaddb <= "110010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001011";
				elsif cntr ="000001001011" THEN
				      ioadda <= "010010111";
				      ioaddb <= "110010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001100";
				elsif cntr ="000001001100" THEN
				      ioadda <= "010011001";
				      ioaddb <= "110011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001101";
				elsif cntr ="000001001101" THEN
				      ioadda <= "010011011";
				      ioaddb <= "110011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001110";
				elsif cntr ="000001001110" THEN
				      ioadda <= "010011101";
				      ioaddb <= "110011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001001111";
				elsif cntr ="000001001111" THEN
				      ioadda <= "010011111";
				      ioaddb <= "110011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010000";
				elsif cntr ="000001010000" THEN
				      ioadda <= "010100001";
				      ioaddb <= "110100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010001";
				elsif cntr ="000001010001" THEN
				      ioadda <= "010100011";
				      ioaddb <= "110100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010010";
				elsif cntr ="000001010010" THEN
				      ioadda <= "010100101";
				      ioaddb <= "110100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010011";
				elsif cntr ="000001010011" THEN
				      ioadda <= "010100111";
				      ioaddb <= "110100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010100";
				elsif cntr ="000001010100" THEN
				      ioadda <= "010101001";
				      ioaddb <= "110101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010101";
				elsif cntr ="000001010101" THEN
				      ioadda <= "010101011";
				      ioaddb <= "110101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010110";
				elsif cntr ="000001010110" THEN
				      ioadda <= "010101101";
				      ioaddb <= "110101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001010111";
				elsif cntr ="000001010111" THEN
				      ioadda <= "010101111";
				      ioaddb <= "110101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011000";
				elsif cntr ="000001011000" THEN
				      ioadda <= "010110001";
				      ioaddb <= "110110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011001";
				elsif cntr ="000001011001" THEN
				      ioadda <= "010110011";
				      ioaddb <= "110110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011010";
				elsif cntr ="000001011010" THEN
				      ioadda <= "010110101";
				      ioaddb <= "110110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011011";
				elsif cntr ="000001011011" THEN
				      ioadda <= "010110111";
				      ioaddb <= "110110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011100";
				elsif cntr ="000001011100" THEN
				      ioadda <= "010111001";
				      ioaddb <= "110111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011101";
				elsif cntr ="000001011101" THEN
				      ioadda <= "010111011";
				      ioaddb <= "110111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011110";
				elsif cntr ="000001011110" THEN
				      ioadda <= "010111101";
				      ioaddb <= "110111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001011111";
				elsif cntr ="000001011111" THEN
				      ioadda <= "010111111";
				      ioaddb <= "110111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100000";
				elsif cntr ="000001100000" THEN
				      ioadda <= "011000001";
				      ioaddb <= "111000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100001";
				elsif cntr ="000001100001" THEN
				      ioadda <= "011000011";
				      ioaddb <= "111000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100010";
				elsif cntr ="000001100010" THEN
				      ioadda <= "011000101";
				      ioaddb <= "111000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100011";
				elsif cntr ="000001100011" THEN
				      ioadda <= "011000111";
				      ioaddb <= "111000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100100";
				elsif cntr ="000001100100" THEN
				      ioadda <= "011001001";
				      ioaddb <= "111001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100101";
				elsif cntr ="000001100101" THEN
				      ioadda <= "011001011";
				      ioaddb <= "111001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100110";
				elsif cntr ="000001100110" THEN
				      ioadda <= "011001101";
				      ioaddb <= "111001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001100111";
				elsif cntr ="000001100111" THEN
				      ioadda <= "011001111";
				      ioaddb <= "111001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101000";
				elsif cntr ="000001101000" THEN
				      ioadda <= "011010001";
				      ioaddb <= "111010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101001";
				elsif cntr ="000001101001" THEN
				      ioadda <= "011010011";
				      ioaddb <= "111010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101010";
				elsif cntr ="000001101010" THEN
				      ioadda <= "011010101";
				      ioaddb <= "111010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101011";
				elsif cntr ="000001101011" THEN
				      ioadda <= "011010111";
				      ioaddb <= "111010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101100";
				elsif cntr ="000001101100" THEN
				      ioadda <= "011011001";
				      ioaddb <= "111011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101101";
				elsif cntr ="000001101101" THEN
				      ioadda <= "011011011";
				      ioaddb <= "111011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101110";
				elsif cntr ="000001101110" THEN
				      ioadda <= "011011101";
				      ioaddb <= "111011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001101111";
				elsif cntr ="000001101111" THEN
				      ioadda <= "011011111";
				      ioaddb <= "111011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110000";
				elsif cntr ="000001110000" THEN
				      ioadda <= "011100001";
				      ioaddb <= "111100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110001";
				elsif cntr ="000001110001" THEN
				      ioadda <= "011100011";
				      ioaddb <= "111100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110010";
				elsif cntr ="000001110010" THEN
				      ioadda <= "011100101";
				      ioaddb <= "111100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110011";
				elsif cntr ="000001110011" THEN
				      ioadda <= "011100111";
				      ioaddb <= "111100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110100";
				elsif cntr ="000001110100" THEN
				      ioadda <= "011101001";
				      ioaddb <= "111101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110101";
				elsif cntr ="000001110101" THEN
				      ioadda <= "011101011";
				      ioaddb <= "111101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110110";
				elsif cntr ="000001110110" THEN
				      ioadda <= "011101101";
				      ioaddb <= "111101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001110111";
				elsif cntr ="000001110111" THEN
				      ioadda <= "011101111";
				      ioaddb <= "111101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111000";
				elsif cntr ="000001111000" THEN
				      ioadda <= "011110001";
				      ioaddb <= "111110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111001";
				elsif cntr ="000001111001" THEN
				      ioadda <= "011110011";
				      ioaddb <= "111110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111010";
				elsif cntr ="000001111010" THEN
				      ioadda <= "011110101";
				      ioaddb <= "111110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111011";
				elsif cntr ="000001111011" THEN
				      ioadda <= "011110111";
				      ioaddb <= "111110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111100";
				elsif cntr ="000001111100" THEN
				      ioadda <= "011111001";
				      ioaddb <= "111111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111101";
				elsif cntr ="000001111101" THEN
				      ioadda <= "011111011";
				      ioaddb <= "111111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111110";
				elsif cntr ="000001111110" THEN
				      ioadda <= "011111101";
				      ioaddb <= "111111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000001111111";
				elsif cntr ="000001111111" THEN
				      ioadda <= "011111111";
				      ioaddb <= "111111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010000000";
				elsif cntr ="000010000000" THEN			
				      ioadda <= "000000000";      
				      ioaddb <= "100000000";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010000001";
				elsif cntr ="000010000001" THEN			
				      ioadda <= "000000010";      
				      ioaddb <= "100000010";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010000010";
				elsif cntr ="000010000010" THEN		
				      ioadda <= "000000100";      
				      ioaddb <= "100000100";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000010000011";      
				elsif cntr ="000010000011" THEN		      
				      ioadda <= "000000110";      
				      ioaddb <= "100000110";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000010000100";            
				elsif cntr ="000010000100" THEN		        
				      ioadda <= "000001000";      
				      ioaddb <= "100001000";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000010000101";             
				elsif cntr ="000010000101" THEN		      
				      ioadda <= "000001010";      
				      ioaddb <= "100001010";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "000010000110";             
				elsif cntr ="000010000110" THEN		      
				      ioadda <= "000001100";      
				      ioaddb <= "100001100";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000010000111";                  
				elsif cntr ="000010000111" THEN		           
				      ioadda <= "000001110";      
				      ioaddb <= "100001110";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000010001000";       
				elsif cntr ="000010001000" THEN		
				      ioadda <= "000010000";
				      ioaddb <= "100010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				      
				      
				      
				      cntr <= "000010001001";
				elsif cntr ="000010001001" THEN
				      ioadda <= "000010010";
				      ioaddb <= "100010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001010";
				elsif cntr ="000010001010" THEN
				      ioadda <= "000010100";
				      ioaddb <= "100010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001011";
				elsif cntr ="000010001011" THEN
				      ioadda <= "000010110";
				      ioaddb <= "100010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001100";
				elsif cntr ="000010001100" THEN
				      ioadda <= "000011000";
				      ioaddb <= "100011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001101";
				elsif cntr ="000010001101" THEN
				      ioadda <= "000011010";
				      ioaddb <= "100011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001110";
				elsif cntr ="000010001110" THEN
				      ioadda <= "000011100";
				      ioaddb <= "100011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010001111";
				elsif cntr ="000010001111" THEN
				      ioadda <= "000011110";
				      ioaddb <= "100011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010000";
				elsif cntr ="000010010000" THEN
				      ioadda <= "000100000";
				      ioaddb <= "100100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010001";
				elsif cntr ="000010010001" THEN
				      ioadda <= "000100010";
				      ioaddb <= "100100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010010";
				elsif cntr ="000010010010" THEN
				      ioadda <= "000100100";
				      ioaddb <= "100100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010011";
				elsif cntr ="000010010011" THEN
				      ioadda <= "000100110";
				      ioaddb <= "100100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010100";
				elsif cntr ="000010010100" THEN
				      ioadda <= "000101000";
				      ioaddb <= "100101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010101";
				elsif cntr ="000010010101" THEN
				      ioadda <= "000101010";
				      ioaddb <= "100101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010110";
				elsif cntr ="000010010110" THEN
				      ioadda <= "000101100";
				      ioaddb <= "100101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010010111";
				elsif cntr ="000010010111" THEN
				      ioadda <= "000101110";
				      ioaddb <= "100101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011000";
				elsif cntr ="000010011000" THEN
				      ioadda <= "000110000";
				      ioaddb <= "100110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011001";
				elsif cntr ="000010011001" THEN
				      ioadda <= "000110010";
				      ioaddb <= "100110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011010";
				elsif cntr ="000010011010" THEN
				      ioadda <= "000110100";
				      ioaddb <= "100110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011011";
				elsif cntr ="000010011011" THEN
				      ioadda <= "000110110";
				      ioaddb <= "100110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011100";
				elsif cntr ="000010011100" THEN
				      ioadda <= "000111000";
				      ioaddb <= "100111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011101";
				elsif cntr ="000010011101" THEN
				      ioadda <= "000111010";
				      ioaddb <= "100111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011110";
				elsif cntr ="000010011110" THEN
				      ioadda <= "000111100";
				      ioaddb <= "100111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010011111";
				elsif cntr ="000010011111" THEN
				      ioadda <= "000111110";
				      ioaddb <= "100111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100000";
				elsif cntr ="000010100000" THEN
				      ioadda <= "001000000";
				      ioaddb <= "101000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100001";
				elsif cntr ="000010100001" THEN
				      ioadda <= "001000010";
				      ioaddb <= "101000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100010";
				elsif cntr ="000010100010" THEN
				      ioadda <= "001000100";
				      ioaddb <= "101000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100011";
				elsif cntr ="000010100011" THEN
				      ioadda <= "001000110";
				      ioaddb <= "101000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100100";
				elsif cntr ="000010100100" THEN
				      ioadda <= "001001000";
				      ioaddb <= "101001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100101";
				elsif cntr ="000010100101" THEN
				      ioadda <= "001001010";
				      ioaddb <= "101001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100110";
				elsif cntr ="000010100110" THEN
				      ioadda <= "001001100";
				      ioaddb <= "101001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010100111";
				elsif cntr ="000010100111" THEN
				      ioadda <= "001001110";
				      ioaddb <= "101001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101000";
				elsif cntr ="000010101000" THEN
				      ioadda <= "001010000";
				      ioaddb <= "101010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101001";
				elsif cntr ="000010101001" THEN
				      ioadda <= "001010010";
				      ioaddb <= "101010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101010";
				elsif cntr ="000010101010" THEN
				      ioadda <= "001010100";
				      ioaddb <= "101010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101011";
				elsif cntr ="000010101011" THEN
				      ioadda <= "001010110";
				      ioaddb <= "101010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101100";
				elsif cntr ="000010101100" THEN
				      ioadda <= "001011000";
				      ioaddb <= "101011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101101";
				elsif cntr ="000010101101" THEN
				      ioadda <= "001011010";
				      ioaddb <= "101011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101110";
				elsif cntr ="000010101110" THEN
				      ioadda <= "001011100";
				      ioaddb <= "101011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010101111";
				elsif cntr ="000010101111" THEN
				      ioadda <= "001011110";
				      ioaddb <= "101011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110000";
				elsif cntr ="000010110000" THEN
				      ioadda <= "001100000";
				      ioaddb <= "101100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110001";
				elsif cntr ="000010110001" THEN
				      ioadda <= "001100010";
				      ioaddb <= "101100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110010";
				elsif cntr ="000010110010" THEN
				      ioadda <= "001100100";
				      ioaddb <= "101100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110011";
				elsif cntr ="000010110011" THEN
				      ioadda <= "001100110";
				      ioaddb <= "101100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110100";
				elsif cntr ="000010110100" THEN
				      ioadda <= "001101000";
				      ioaddb <= "101101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110101";
				elsif cntr ="000010110101" THEN
				      ioadda <= "001101010";
				      ioaddb <= "101101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110110";
				elsif cntr ="000010110110" THEN
				      ioadda <= "001101100";
				      ioaddb <= "101101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010110111";
				elsif cntr ="000010110111" THEN
				      ioadda <= "001101110";
				      ioaddb <= "101101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111000";
				elsif cntr ="000010111000" THEN
				      ioadda <= "001110000";
				      ioaddb <= "101110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111001";
				elsif cntr ="000010111001" THEN
				      ioadda <= "001110010";
				      ioaddb <= "101110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111010";
				elsif cntr ="000010111010" THEN
				      ioadda <= "001110100";
				      ioaddb <= "101110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111011";
				elsif cntr ="000010111011" THEN
				      ioadda <= "001110110";
				      ioaddb <= "101110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111100";
				elsif cntr ="000010111100" THEN
				      ioadda <= "001111000";
				      ioaddb <= "101111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111101";
				elsif cntr ="000010111101" THEN
				      ioadda <= "001111010";
				      ioaddb <= "101111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111110";
				elsif cntr ="000010111110" THEN
				      ioadda <= "001111100";
				      ioaddb <= "101111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000010111111";
				elsif cntr ="000010111111" THEN
				      ioadda <= "001111110";
				      ioaddb <= "101111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000000";
				elsif cntr ="000011000000" THEN
				      ioadda <= "010000000";
				      ioaddb <= "110000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000001";
				elsif cntr ="000011000001" THEN
				      ioadda <= "010000010";
				      ioaddb <= "110000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000010";
				elsif cntr ="000011000010" THEN
				      ioadda <= "010000100";
				      ioaddb <= "110000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000011";
				elsif cntr ="000011000011" THEN
				      ioadda <= "010000110";
				      ioaddb <= "110000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000100";
				elsif cntr ="000011000100" THEN
				      ioadda <= "010001000";
				      ioaddb <= "110001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000101";
				elsif cntr ="000011000101" THEN
				      ioadda <= "010001010";
				      ioaddb <= "110001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000110";
				elsif cntr ="000011000110" THEN
				      ioadda <= "010001100";
				      ioaddb <= "110001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011000111";
				elsif cntr ="000011000111" THEN
				      ioadda <= "010001110";
				      ioaddb <= "110001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001000";
				elsif cntr ="000011001000" THEN
				      ioadda <= "010010000";
				      ioaddb <= "110010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001001";
				elsif cntr ="000011001001" THEN
				      ioadda <= "010010010";
				      ioaddb <= "110010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001010";
				elsif cntr ="000011001010" THEN
				      ioadda <= "010010100";
				      ioaddb <= "110010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001011";
				elsif cntr ="000011001011" THEN
				      ioadda <= "010010110";
				      ioaddb <= "110010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001100";
				elsif cntr ="000011001100" THEN
				      ioadda <= "010011000";
				      ioaddb <= "110011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001101";
				elsif cntr ="000011001101" THEN
				      ioadda <= "010011010";
				      ioaddb <= "110011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001110";
				elsif cntr ="000011001110" THEN
				      ioadda <= "010011100";
				      ioaddb <= "110011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011001111";
				elsif cntr ="000011001111" THEN
				      ioadda <= "010011110";
				      ioaddb <= "110011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010000";
				elsif cntr ="000011010000" THEN
				      ioadda <= "010100000";
				      ioaddb <= "110100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010001";
				elsif cntr ="000011010001" THEN
				      ioadda <= "010100010";
				      ioaddb <= "110100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010010";
				elsif cntr ="000011010010" THEN
				      ioadda <= "010100100";
				      ioaddb <= "110100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010011";
				elsif cntr ="000011010011" THEN
				      ioadda <= "010100110";
				      ioaddb <= "110100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010100";
				elsif cntr ="000011010100" THEN
				      ioadda <= "010101000";
				      ioaddb <= "110101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010101";
				elsif cntr ="000011010101" THEN
				      ioadda <= "010101010";
				      ioaddb <= "110101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010110";
				elsif cntr ="000011010110" THEN
				      ioadda <= "010101100";
				      ioaddb <= "110101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011010111";
				elsif cntr ="000011010111" THEN
				      ioadda <= "010101110";
				      ioaddb <= "110101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011000";
				elsif cntr ="000011011000" THEN
				      ioadda <= "010110000";
				      ioaddb <= "110110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011001";
				elsif cntr ="000011011001" THEN
				      ioadda <= "010110010";
				      ioaddb <= "110110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011010";
				elsif cntr ="000011011010" THEN
				      ioadda <= "010110100";
				      ioaddb <= "110110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011011";
				elsif cntr ="000011011011" THEN
				      ioadda <= "010110110";
				      ioaddb <= "110110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011100";
				elsif cntr ="000011011100" THEN
				      ioadda <= "010111000";
				      ioaddb <= "110111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011101";
				elsif cntr ="000011011101" THEN
				      ioadda <= "010111010";
				      ioaddb <= "110111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011110";
				elsif cntr ="000011011110" THEN
				      ioadda <= "010111100";
				      ioaddb <= "110111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011011111";
				elsif cntr ="000011011111" THEN
				      ioadda <= "010111110";
				      ioaddb <= "110111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100000";
				elsif cntr ="000011100000" THEN
				      ioadda <= "011000000";
				      ioaddb <= "111000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100001";
				elsif cntr ="000011100001" THEN
				      ioadda <= "011000010";
				      ioaddb <= "111000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100010";
				elsif cntr ="000011100010" THEN
				      ioadda <= "011000100";
				      ioaddb <= "111000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100011";
				elsif cntr ="000011100011" THEN
				      ioadda <= "011000110";
				      ioaddb <= "111000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100100";
				elsif cntr ="000011100100" THEN
				      ioadda <= "011001000";
				      ioaddb <= "111001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100101";
				elsif cntr ="000011100101" THEN
				      ioadda <= "011001010";
				      ioaddb <= "111001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100110";
				elsif cntr ="000011100110" THEN
				      ioadda <= "011001100";
				      ioaddb <= "111001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011100111";
				elsif cntr ="000011100111" THEN
				      ioadda <= "011001110";
				      ioaddb <= "111001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101000";
				elsif cntr ="000011101000" THEN
				      ioadda <= "011010000";
				      ioaddb <= "111010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101001";
				elsif cntr ="000011101001" THEN
				      ioadda <= "011010010";
				      ioaddb <= "111010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101010";
				elsif cntr ="000011101010" THEN
				      ioadda <= "011010100";
				      ioaddb <= "111010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101011";
				elsif cntr ="000011101011" THEN
				      ioadda <= "011010110";
				      ioaddb <= "111010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101100";
				elsif cntr ="000011101100" THEN
				      ioadda <= "011011000";
				      ioaddb <= "111011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101101";
				elsif cntr ="000011101101" THEN
				      ioadda <= "011011010";
				      ioaddb <= "111011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101110";
				elsif cntr ="000011101110" THEN
				      ioadda <= "011011100";
				      ioaddb <= "111011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011101111";
				elsif cntr ="000011101111" THEN
				      ioadda <= "011011110";
				      ioaddb <= "111011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110000";
				elsif cntr ="000011110000" THEN
				      ioadda <= "011100000";
				      ioaddb <= "111100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110001";
				elsif cntr ="000011110001" THEN
				      ioadda <= "011100010";
				      ioaddb <= "111100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110010";
				elsif cntr ="000011110010" THEN
				      ioadda <= "011100100";
				      ioaddb <= "111100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110011";
				elsif cntr ="000011110011" THEN
				      ioadda <= "011100110";
				      ioaddb <= "111100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110100";
				elsif cntr ="000011110100" THEN
				      ioadda <= "011101000";
				      ioaddb <= "111101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110101";
				elsif cntr ="000011110101" THEN
				      ioadda <= "011101010";
				      ioaddb <= "111101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110110";
				elsif cntr ="000011110110" THEN
				      ioadda <= "011101100";
				      ioaddb <= "111101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011110111";
				elsif cntr ="000011110111" THEN
				      ioadda <= "011101110";
				      ioaddb <= "111101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111000";
				elsif cntr ="000011111000" THEN
				      ioadda <= "011110000";
				      ioaddb <= "111110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111001";
				elsif cntr ="000011111001" THEN
				      ioadda <= "011110010";
				      ioaddb <= "111110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111010";
				elsif cntr ="000011111010" THEN
				      ioadda <= "011110100";
				      ioaddb <= "111110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111011";
				elsif cntr ="000011111011" THEN
				      ioadda <= "011110110";
				      ioaddb <= "111110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111100";
				elsif cntr ="000011111100" THEN
				      ioadda <= "011111000";
				      ioaddb <= "111111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111101";
				elsif cntr ="000011111101" THEN
				      ioadda <= "011111010";
				      ioaddb <= "111111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111110";
				elsif cntr ="000011111110" THEN
				      ioadda <= "011111100";
				      ioaddb <= "111111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000011111111";
				elsif cntr ="000011111111" THEN
				      ioadda <= "011111110";
				      ioaddb <= "111111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100000000";
				elsif cntr ="000100000000" THEN														
				      ioadda <= "000000000";      
				      ioaddb <= "100000001";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100000001";
				elsif cntr ="000100000001" THEN	
				      ioadda <= "000000010";      
				      ioaddb <= "100000011";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100000010";
				elsif cntr ="000100000010" THEN	
				      ioadda <= "000000100";      
				      ioaddb <= "100000101";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000100000011";      
				elsif cntr ="000100000011" THEN	      
				      ioadda <= "000000110";      
				      ioaddb <= "100000111";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000100000100";            
				elsif cntr ="000100000100" THEN	         
				      ioadda <= "000001000";      
				      ioaddb <= "100001001";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000100000101";               
				elsif cntr ="000100000101" THEN	            
				      ioadda <= "000001010";      
				      ioaddb <= "100001011";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "000100000110";                
				elsif cntr ="000100000110" THEN	             
				      ioadda <= "000001100";      
				      ioaddb <= "100001101";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000100000111";          
				elsif cntr ="000100000111" THEN	       
				      ioadda <= "000001110";      
				      ioaddb <= "100001111";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                   
				                                   
				                                   
				      cntr <= "000100001000";      
				elsif cntr ="000100001000" THEN	   
				      ioadda <= "000010000";
				      ioaddb <= "100010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				      
				      
				      
				      cntr <= "000100001001";
				elsif cntr ="000100001001" THEN
				      ioadda <= "000010010";
				      ioaddb <= "100010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001010";
				elsif cntr ="000100001010" THEN
				      ioadda <= "000010100";
				      ioaddb <= "100010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001011";
				elsif cntr ="000100001011" THEN
				      ioadda <= "000010110";
				      ioaddb <= "100010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001100";
				elsif cntr ="000100001100" THEN
				      ioadda <= "000011000";
				      ioaddb <= "100011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001101";
				elsif cntr ="000100001101" THEN
				      ioadda <= "000011010";
				      ioaddb <= "100011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001110";
				elsif cntr ="000100001110" THEN
				      ioadda <= "000011100";
				      ioaddb <= "100011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100001111";
				elsif cntr ="000100001111" THEN
				      ioadda <= "000011110";
				      ioaddb <= "100011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010000";
				elsif cntr ="000100010000" THEN
				      ioadda <= "000100000";
				      ioaddb <= "100100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010001";
				elsif cntr ="000100010001" THEN
				      ioadda <= "000100010";
				      ioaddb <= "100100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010010";
				elsif cntr ="000100010010" THEN
				      ioadda <= "000100100";
				      ioaddb <= "100100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010011";
				elsif cntr ="000100010011" THEN
				      ioadda <= "000100110";
				      ioaddb <= "100100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010100";
				elsif cntr ="000100010100" THEN
				      ioadda <= "000101000";
				      ioaddb <= "100101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010101";
				elsif cntr ="000100010101" THEN
				      ioadda <= "000101010";
				      ioaddb <= "100101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010110";
				elsif cntr ="000100010110" THEN
				      ioadda <= "000101100";
				      ioaddb <= "100101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100010111";
				elsif cntr ="000100010111" THEN
				      ioadda <= "000101110";
				      ioaddb <= "100101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011000";
				elsif cntr ="000100011000" THEN
				      ioadda <= "000110000";
				      ioaddb <= "100110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011001";
				elsif cntr ="000100011001" THEN
				      ioadda <= "000110010";
				      ioaddb <= "100110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011010";
				elsif cntr ="000100011010" THEN
				      ioadda <= "000110100";
				      ioaddb <= "100110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011011";
				elsif cntr ="000100011011" THEN
				      ioadda <= "000110110";
				      ioaddb <= "100110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011100";
				elsif cntr ="000100011100" THEN
				      ioadda <= "000111000";
				      ioaddb <= "100111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011101";
				elsif cntr ="000100011101" THEN
				      ioadda <= "000111010";
				      ioaddb <= "100111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011110";
				elsif cntr ="000100011110" THEN
				      ioadda <= "000111100";
				      ioaddb <= "100111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100011111";
				elsif cntr ="000100011111" THEN
				      ioadda <= "000111110";
				      ioaddb <= "100111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100000";
				elsif cntr ="000100100000" THEN
				      ioadda <= "001000000";
				      ioaddb <= "101000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100001";
				elsif cntr ="000100100001" THEN
				      ioadda <= "001000010";
				      ioaddb <= "101000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100010";
				elsif cntr ="000100100010" THEN
				      ioadda <= "001000100";
				      ioaddb <= "101000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100011";
				elsif cntr ="000100100011" THEN
				      ioadda <= "001000110";
				      ioaddb <= "101000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100100";
				elsif cntr ="000100100100" THEN
				      ioadda <= "001001000";
				      ioaddb <= "101001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100101";
				elsif cntr ="000100100101" THEN
				      ioadda <= "001001010";
				      ioaddb <= "101001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100110";
				elsif cntr ="000100100110" THEN
				      ioadda <= "001001100";
				      ioaddb <= "101001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100100111";
				elsif cntr ="000100100111" THEN
				      ioadda <= "001001110";
				      ioaddb <= "101001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101000";
				elsif cntr ="000100101000" THEN
				      ioadda <= "001010000";
				      ioaddb <= "101010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101001";
				elsif cntr ="000100101001" THEN
				      ioadda <= "001010010";
				      ioaddb <= "101010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101010";
				elsif cntr ="000100101010" THEN
				      ioadda <= "001010100";
				      ioaddb <= "101010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101011";
				elsif cntr ="000100101011" THEN
				      ioadda <= "001010110";
				      ioaddb <= "101010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101100";
				elsif cntr ="000100101100" THEN
				      ioadda <= "001011000";
				      ioaddb <= "101011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101101";
				elsif cntr ="000100101101" THEN
				      ioadda <= "001011010";
				      ioaddb <= "101011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101110";
				elsif cntr ="000100101110" THEN
				      ioadda <= "001011100";
				      ioaddb <= "101011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100101111";
				elsif cntr ="000100101111" THEN
				      ioadda <= "001011110";
				      ioaddb <= "101011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110000";
				elsif cntr ="000100110000" THEN
				      ioadda <= "001100000";
				      ioaddb <= "101100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110001";
				elsif cntr ="000100110001" THEN
				      ioadda <= "001100010";
				      ioaddb <= "101100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110010";
				elsif cntr ="000100110010" THEN
				      ioadda <= "001100100";
				      ioaddb <= "101100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110011";
				elsif cntr ="000100110011" THEN
				      ioadda <= "001100110";
				      ioaddb <= "101100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110100";
				elsif cntr ="000100110100" THEN
				      ioadda <= "001101000";
				      ioaddb <= "101101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110101";
				elsif cntr ="000100110101" THEN
				      ioadda <= "001101010";
				      ioaddb <= "101101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110110";
				elsif cntr ="000100110110" THEN
				      ioadda <= "001101100";
				      ioaddb <= "101101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100110111";
				elsif cntr ="000100110111" THEN
				      ioadda <= "001101110";
				      ioaddb <= "101101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111000";
				elsif cntr ="000100111000" THEN
				      ioadda <= "001110000";
				      ioaddb <= "101110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111001";
				elsif cntr ="000100111001" THEN
				      ioadda <= "001110010";
				      ioaddb <= "101110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111010";
				elsif cntr ="000100111010" THEN
				      ioadda <= "001110100";
				      ioaddb <= "101110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111011";
				elsif cntr ="000100111011" THEN
				      ioadda <= "001110110";
				      ioaddb <= "101110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111100";
				elsif cntr ="000100111100" THEN
				      ioadda <= "001111000";
				      ioaddb <= "101111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111101";
				elsif cntr ="000100111101" THEN
				      ioadda <= "001111010";
				      ioaddb <= "101111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111110";
				elsif cntr ="000100111110" THEN
				      ioadda <= "001111100";
				      ioaddb <= "101111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000100111111";
				elsif cntr ="000100111111" THEN
				      ioadda <= "001111110";
				      ioaddb <= "101111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000000";
				elsif cntr ="000101000000" THEN
				      ioadda <= "010000000";
				      ioaddb <= "110000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000001";
				elsif cntr ="000101000001" THEN
				      ioadda <= "010000010";
				      ioaddb <= "110000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000010";
				elsif cntr ="000101000010" THEN
				      ioadda <= "010000100";
				      ioaddb <= "110000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000011";
				elsif cntr ="000101000011" THEN
				      ioadda <= "010000110";
				      ioaddb <= "110000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000100";
				elsif cntr ="000101000100" THEN
				      ioadda <= "010001000";
				      ioaddb <= "110001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000101";
				elsif cntr ="000101000101" THEN
				      ioadda <= "010001010";
				      ioaddb <= "110001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000110";
				elsif cntr ="000101000110" THEN
				      ioadda <= "010001100";
				      ioaddb <= "110001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101000111";
				elsif cntr ="000101000111" THEN
				      ioadda <= "010001110";
				      ioaddb <= "110001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001000";
				elsif cntr ="000101001000" THEN
				      ioadda <= "010010000";
				      ioaddb <= "110010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001001";
				elsif cntr ="000101001001" THEN
				      ioadda <= "010010010";
				      ioaddb <= "110010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001010";
				elsif cntr ="000101001010" THEN
				      ioadda <= "010010100";
				      ioaddb <= "110010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001011";
				elsif cntr ="000101001011" THEN
				      ioadda <= "010010110";
				      ioaddb <= "110010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001100";
				elsif cntr ="000101001100" THEN
				      ioadda <= "010011000";
				      ioaddb <= "110011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001101";
				elsif cntr ="000101001101" THEN
				      ioadda <= "010011010";
				      ioaddb <= "110011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001110";
				elsif cntr ="000101001110" THEN
				      ioadda <= "010011100";
				      ioaddb <= "110011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101001111";
				elsif cntr ="000101001111" THEN
				      ioadda <= "010011110";
				      ioaddb <= "110011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010000";
				elsif cntr ="000101010000" THEN
				      ioadda <= "010100000";
				      ioaddb <= "110100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010001";
				elsif cntr ="000101010001" THEN
				      ioadda <= "010100010";
				      ioaddb <= "110100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010010";
				elsif cntr ="000101010010" THEN
				      ioadda <= "010100100";
				      ioaddb <= "110100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010011";
				elsif cntr ="000101010011" THEN
				      ioadda <= "010100110";
				      ioaddb <= "110100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010100";
				elsif cntr ="000101010100" THEN
				      ioadda <= "010101000";
				      ioaddb <= "110101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010101";
				elsif cntr ="000101010101" THEN
				      ioadda <= "010101010";
				      ioaddb <= "110101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010110";
				elsif cntr ="000101010110" THEN
				      ioadda <= "010101100";
				      ioaddb <= "110101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101010111";
				elsif cntr ="000101010111" THEN
				      ioadda <= "010101110";
				      ioaddb <= "110101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011000";
				elsif cntr ="000101011000" THEN
				      ioadda <= "010110000";
				      ioaddb <= "110110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011001";
				elsif cntr ="000101011001" THEN
				      ioadda <= "010110010";
				      ioaddb <= "110110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011010";
				elsif cntr ="000101011010" THEN
				      ioadda <= "010110100";
				      ioaddb <= "110110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011011";
				elsif cntr ="000101011011" THEN
				      ioadda <= "010110110";
				      ioaddb <= "110110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011100";
				elsif cntr ="000101011100" THEN
				      ioadda <= "010111000";
				      ioaddb <= "110111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011101";
				elsif cntr ="000101011101" THEN
				      ioadda <= "010111010";
				      ioaddb <= "110111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011110";
				elsif cntr ="000101011110" THEN
				      ioadda <= "010111100";
				      ioaddb <= "110111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101011111";
				elsif cntr ="000101011111" THEN
				      ioadda <= "010111110";
				      ioaddb <= "110111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100000";
				elsif cntr ="000101100000" THEN
				      ioadda <= "011000000";
				      ioaddb <= "111000001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100001";
				elsif cntr ="000101100001" THEN
				      ioadda <= "011000010";
				      ioaddb <= "111000011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100010";
				elsif cntr ="000101100010" THEN
				      ioadda <= "011000100";
				      ioaddb <= "111000101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100011";
				elsif cntr ="000101100011" THEN
				      ioadda <= "011000110";
				      ioaddb <= "111000111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100100";
				elsif cntr ="000101100100" THEN
				      ioadda <= "011001000";
				      ioaddb <= "111001001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100101";
				elsif cntr ="000101100101" THEN
				      ioadda <= "011001010";
				      ioaddb <= "111001011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100110";
				elsif cntr ="000101100110" THEN
				      ioadda <= "011001100";
				      ioaddb <= "111001101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101100111";
				elsif cntr ="000101100111" THEN
				      ioadda <= "011001110";
				      ioaddb <= "111001111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101000";
				elsif cntr ="000101101000" THEN
				      ioadda <= "011010000";
				      ioaddb <= "111010001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101001";
				elsif cntr ="000101101001" THEN
				      ioadda <= "011010010";
				      ioaddb <= "111010011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101010";
				elsif cntr ="000101101010" THEN
				      ioadda <= "011010100";
				      ioaddb <= "111010101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101011";
				elsif cntr ="000101101011" THEN
				      ioadda <= "011010110";
				      ioaddb <= "111010111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101100";
				elsif cntr ="000101101100" THEN
				      ioadda <= "011011000";
				      ioaddb <= "111011001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101101";
				elsif cntr ="000101101101" THEN
				      ioadda <= "011011010";
				      ioaddb <= "111011011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101110";
				elsif cntr ="000101101110" THEN
				      ioadda <= "011011100";
				      ioaddb <= "111011101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101101111";
				elsif cntr ="000101101111" THEN
				      ioadda <= "011011110";
				      ioaddb <= "111011111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110000";
				elsif cntr ="000101110000" THEN
				      ioadda <= "011100000";
				      ioaddb <= "111100001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110001";
				elsif cntr ="000101110001" THEN
				      ioadda <= "011100010";
				      ioaddb <= "111100011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110010";
				elsif cntr ="000101110010" THEN
				      ioadda <= "011100100";
				      ioaddb <= "111100101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110011";
				elsif cntr ="000101110011" THEN
				      ioadda <= "011100110";
				      ioaddb <= "111100111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110100";
				elsif cntr ="000101110100" THEN
				      ioadda <= "011101000";
				      ioaddb <= "111101001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110101";
				elsif cntr ="000101110101" THEN
				      ioadda <= "011101010";
				      ioaddb <= "111101011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110110";
				elsif cntr ="000101110110" THEN
				      ioadda <= "011101100";
				      ioaddb <= "111101101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101110111";
				elsif cntr ="000101110111" THEN
				      ioadda <= "011101110";
				      ioaddb <= "111101111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111000";
				elsif cntr ="000101111000" THEN
				      ioadda <= "011110000";
				      ioaddb <= "111110001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111001";
				elsif cntr ="000101111001" THEN
				      ioadda <= "011110010";
				      ioaddb <= "111110011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111010";
				elsif cntr ="000101111010" THEN
				      ioadda <= "011110100";
				      ioaddb <= "111110101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111011";
				elsif cntr ="000101111011" THEN
				      ioadda <= "011110110";
				      ioaddb <= "111110111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111100";
				elsif cntr ="000101111100" THEN
				      ioadda <= "011111000";
				      ioaddb <= "111111001";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111101";
				elsif cntr ="000101111101" THEN
				      ioadda <= "011111010";
				      ioaddb <= "111111011";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111110";
				elsif cntr ="000101111110" THEN
				      ioadda <= "011111100";
				      ioaddb <= "111111101";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000101111111";
				elsif cntr ="000101111111" THEN
				      ioadda <= "011111110";
				      ioaddb <= "111111111";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110000000";
				elsif cntr ="000110000000" THEN													
				      ioadda <= "000000001";      
				      ioaddb <= "100000000";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110000001";
				elsif cntr ="000110000001" THEN		
				      ioadda <= "000000011";      
				      ioaddb <= "100000010";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110000010";
				elsif cntr ="000110000010" THEN		
				      ioadda <= "000000101";      
				      ioaddb <= "100000100";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				            
				            
				            
				      cntr <= "000110000011";      
				elsif cntr ="000110000011" THEN		      
				      ioadda <= "000000111";      
				      ioaddb <= "100000110";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "000110000100";            
				elsif cntr ="000110000100" THEN		      
				      ioadda <= "000001001";      
				      ioaddb <= "100001000";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "000110000101";              
				elsif cntr ="000110000101" THEN		       
				      ioadda <= "000001011";      
				      ioaddb <= "100001010";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "000110000110";             
				elsif cntr ="000110000110" THEN		      
				      ioadda <= "000001101";      
				      ioaddb <= "100001100";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "000110000111";         
				elsif cntr ="000110000111" THEN	      
				      ioadda <= "000001111";      
				      ioaddb <= "100001110";      
				      bfrjin   <= iodouta;      
				      bfrjplin <= iodoutb;      
				      
				      
				      
				                                   
				                                   
				                                   
				      cntr <= "000110001000";      
				elsif cntr ="000110001000" THEN	   
				      ioadda <= "000010001";
				      ioaddb <= "100010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				
				
				
				      
				      
				      
				      cntr <= "000110001001";
				elsif cntr ="000110001001" THEN
				      ioadda <= "000010011";
				      ioaddb <= "100010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001010";
				elsif cntr ="000110001010" THEN
				      ioadda <= "000010101";
				      ioaddb <= "100010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001011";
				elsif cntr ="000110001011" THEN
				      ioadda <= "000010111";
				      ioaddb <= "100010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001100";
				elsif cntr ="000110001100" THEN
				      ioadda <= "000011001";
				      ioaddb <= "100011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001101";
				elsif cntr ="000110001101" THEN
				      ioadda <= "000011011";
				      ioaddb <= "100011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001110";
				elsif cntr ="000110001110" THEN
				      ioadda <= "000011101";
				      ioaddb <= "100011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110001111";
				elsif cntr ="000110001111" THEN
				      ioadda <= "000011111";
				      ioaddb <= "100011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010000";
				elsif cntr ="000110010000" THEN
				      ioadda <= "000100001";
				      ioaddb <= "100100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010001";
				elsif cntr ="000110010001" THEN
				      ioadda <= "000100011";
				      ioaddb <= "100100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010010";
				elsif cntr ="000110010010" THEN
				      ioadda <= "000100101";
				      ioaddb <= "100100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010011";
				elsif cntr ="000110010011" THEN
				      ioadda <= "000100111";
				      ioaddb <= "100100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010100";
				elsif cntr ="000110010100" THEN
				      ioadda <= "000101001";
				      ioaddb <= "100101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010101";
				elsif cntr ="000110010101" THEN
				      ioadda <= "000101011";
				      ioaddb <= "100101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010110";
				elsif cntr ="000110010110" THEN
				      ioadda <= "000101101";
				      ioaddb <= "100101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110010111";
				elsif cntr ="000110010111" THEN
				      ioadda <= "000101111";
				      ioaddb <= "100101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011000";
				elsif cntr ="000110011000" THEN
				      ioadda <= "000110001";
				      ioaddb <= "100110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011001";
				elsif cntr ="000110011001" THEN
				      ioadda <= "000110011";
				      ioaddb <= "100110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011010";
				elsif cntr ="000110011010" THEN
				      ioadda <= "000110101";
				      ioaddb <= "100110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011011";
				elsif cntr ="000110011011" THEN
				      ioadda <= "000110111";
				      ioaddb <= "100110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011100";
				elsif cntr ="000110011100" THEN
				      ioadda <= "000111001";
				      ioaddb <= "100111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011101";
				elsif cntr ="000110011101" THEN
				      ioadda <= "000111011";
				      ioaddb <= "100111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011110";
				elsif cntr ="000110011110" THEN
				      ioadda <= "000111101";
				      ioaddb <= "100111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110011111";
				elsif cntr ="000110011111" THEN
				      ioadda <= "000111111";
				      ioaddb <= "100111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100000";
				elsif cntr ="000110100000" THEN
				      ioadda <= "001000001";
				      ioaddb <= "101000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100001";
				elsif cntr ="000110100001" THEN
				      ioadda <= "001000011";
				      ioaddb <= "101000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100010";
				elsif cntr ="000110100010" THEN
				      ioadda <= "001000101";
				      ioaddb <= "101000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100011";
				elsif cntr ="000110100011" THEN
				      ioadda <= "001000111";
				      ioaddb <= "101000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100100";
				elsif cntr ="000110100100" THEN
				      ioadda <= "001001001";
				      ioaddb <= "101001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100101";
				elsif cntr ="000110100101" THEN
				      ioadda <= "001001011";
				      ioaddb <= "101001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100110";
				elsif cntr ="000110100110" THEN
				      ioadda <= "001001101";
				      ioaddb <= "101001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110100111";
				elsif cntr ="000110100111" THEN
				      ioadda <= "001001111";
				      ioaddb <= "101001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101000";
				elsif cntr ="000110101000" THEN
				      ioadda <= "001010001";
				      ioaddb <= "101010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101001";
				elsif cntr ="000110101001" THEN
				      ioadda <= "001010011";
				      ioaddb <= "101010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101010";
				elsif cntr ="000110101010" THEN
				      ioadda <= "001010101";
				      ioaddb <= "101010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101011";
				elsif cntr ="000110101011" THEN
				      ioadda <= "001010111";
				      ioaddb <= "101010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101100";
				elsif cntr ="000110101100" THEN
				      ioadda <= "001011001";
				      ioaddb <= "101011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101101";
				elsif cntr ="000110101101" THEN
				      ioadda <= "001011011";
				      ioaddb <= "101011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101110";
				elsif cntr ="000110101110" THEN
				      ioadda <= "001011101";
				      ioaddb <= "101011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110101111";
				elsif cntr ="000110101111" THEN
				      ioadda <= "001011111";
				      ioaddb <= "101011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110000";
				elsif cntr ="000110110000" THEN
				      ioadda <= "001100001";
				      ioaddb <= "101100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110001";
				elsif cntr ="000110110001" THEN
				      ioadda <= "001100011";
				      ioaddb <= "101100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110010";
				elsif cntr ="000110110010" THEN
				      ioadda <= "001100101";
				      ioaddb <= "101100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110011";
				elsif cntr ="000110110011" THEN
				      ioadda <= "001100111";
				      ioaddb <= "101100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110100";
				elsif cntr ="000110110100" THEN
				      ioadda <= "001101001";
				      ioaddb <= "101101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110101";
				elsif cntr ="000110110101" THEN
				      ioadda <= "001101011";
				      ioaddb <= "101101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110110";
				elsif cntr ="000110110110" THEN
				      ioadda <= "001101101";
				      ioaddb <= "101101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110110111";
				elsif cntr ="000110110111" THEN
				      ioadda <= "001101111";
				      ioaddb <= "101101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111000";
				elsif cntr ="000110111000" THEN
				      ioadda <= "001110001";
				      ioaddb <= "101110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111001";
				elsif cntr ="000110111001" THEN
				      ioadda <= "001110011";
				      ioaddb <= "101110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111010";
				elsif cntr ="000110111010" THEN
				      ioadda <= "001110101";
				      ioaddb <= "101110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111011";
				elsif cntr ="000110111011" THEN
				      ioadda <= "001110111";
				      ioaddb <= "101110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111100";
				elsif cntr ="000110111100" THEN
				      ioadda <= "001111001";
				      ioaddb <= "101111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111101";
				elsif cntr ="000110111101" THEN
				      ioadda <= "001111011";
				      ioaddb <= "101111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111110";
				elsif cntr ="000110111110" THEN
				      ioadda <= "001111101";
				      ioaddb <= "101111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000110111111";
				elsif cntr ="000110111111" THEN
				      ioadda <= "001111111";
				      ioaddb <= "101111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000000";
				elsif cntr ="000111000000" THEN
				      ioadda <= "010000001";
				      ioaddb <= "110000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000001";
				elsif cntr ="000111000001" THEN
				      ioadda <= "010000011";
				      ioaddb <= "110000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000010";
				elsif cntr ="000111000010" THEN
				      ioadda <= "010000101";
				      ioaddb <= "110000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000011";
				elsif cntr ="000111000011" THEN
				      ioadda <= "010000111";
				      ioaddb <= "110000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000100";
				elsif cntr ="000111000100" THEN
				      ioadda <= "010001001";
				      ioaddb <= "110001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000101";
				elsif cntr ="000111000101" THEN
				      ioadda <= "010001011";
				      ioaddb <= "110001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000110";
				elsif cntr ="000111000110" THEN
				      ioadda <= "010001101";
				      ioaddb <= "110001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111000111";
				elsif cntr ="000111000111" THEN
				      ioadda <= "010001111";
				      ioaddb <= "110001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001000";
				elsif cntr ="000111001000" THEN
				      ioadda <= "010010001";
				      ioaddb <= "110010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001001";
				elsif cntr ="000111001001" THEN
				      ioadda <= "010010011";
				      ioaddb <= "110010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001010";
				elsif cntr ="000111001010" THEN
				      ioadda <= "010010101";
				      ioaddb <= "110010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001011";
				elsif cntr ="000111001011" THEN
				      ioadda <= "010010111";
				      ioaddb <= "110010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001100";
				elsif cntr ="000111001100" THEN
				      ioadda <= "010011001";
				      ioaddb <= "110011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001101";
				elsif cntr ="000111001101" THEN
				      ioadda <= "010011011";
				      ioaddb <= "110011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001110";
				elsif cntr ="000111001110" THEN
				      ioadda <= "010011101";
				      ioaddb <= "110011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111001111";
				elsif cntr ="000111001111" THEN
				      ioadda <= "010011111";
				      ioaddb <= "110011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010000";
				elsif cntr ="000111010000" THEN
				      ioadda <= "010100001";
				      ioaddb <= "110100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010001";
				elsif cntr ="000111010001" THEN
				      ioadda <= "010100011";
				      ioaddb <= "110100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010010";
				elsif cntr ="000111010010" THEN
				      ioadda <= "010100101";
				      ioaddb <= "110100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010011";
				elsif cntr ="000111010011" THEN
				      ioadda <= "010100111";
				      ioaddb <= "110100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010100";
				elsif cntr ="000111010100" THEN
				      ioadda <= "010101001";
				      ioaddb <= "110101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010101";
				elsif cntr ="000111010101" THEN
				      ioadda <= "010101011";
				      ioaddb <= "110101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010110";
				elsif cntr ="000111010110" THEN
				      ioadda <= "010101101";
				      ioaddb <= "110101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111010111";
				elsif cntr ="000111010111" THEN
				      ioadda <= "010101111";
				      ioaddb <= "110101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011000";
				elsif cntr ="000111011000" THEN
				      ioadda <= "010110001";
				      ioaddb <= "110110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011001";
				elsif cntr ="000111011001" THEN
				      ioadda <= "010110011";
				      ioaddb <= "110110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011010";
				elsif cntr ="000111011010" THEN
				      ioadda <= "010110101";
				      ioaddb <= "110110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011011";
				elsif cntr ="000111011011" THEN
				      ioadda <= "010110111";
				      ioaddb <= "110110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011100";
				elsif cntr ="000111011100" THEN
				      ioadda <= "010111001";
				      ioaddb <= "110111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011101";
				elsif cntr ="000111011101" THEN
				      ioadda <= "010111011";
				      ioaddb <= "110111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011110";
				elsif cntr ="000111011110" THEN
				      ioadda <= "010111101";
				      ioaddb <= "110111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111011111";
				elsif cntr ="000111011111" THEN
				      ioadda <= "010111111";
				      ioaddb <= "110111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100000";
				elsif cntr ="000111100000" THEN
				      ioadda <= "011000001";
				      ioaddb <= "111000000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100001";
				elsif cntr ="000111100001" THEN
				      ioadda <= "011000011";
				      ioaddb <= "111000010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100010";
				elsif cntr ="000111100010" THEN
				      ioadda <= "011000101";
				      ioaddb <= "111000100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100011";
				elsif cntr ="000111100011" THEN
				      ioadda <= "011000111";
				      ioaddb <= "111000110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100100";
				elsif cntr ="000111100100" THEN
				      ioadda <= "011001001";
				      ioaddb <= "111001000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100101";
				elsif cntr ="000111100101" THEN
				      ioadda <= "011001011";
				      ioaddb <= "111001010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100110";
				elsif cntr ="000111100110" THEN
				      ioadda <= "011001101";
				      ioaddb <= "111001100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111100111";
				elsif cntr ="000111100111" THEN
				      ioadda <= "011001111";
				      ioaddb <= "111001110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101000";
				elsif cntr ="000111101000" THEN
				      ioadda <= "011010001";
				      ioaddb <= "111010000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101001";
				elsif cntr ="000111101001" THEN
				      ioadda <= "011010011";
				      ioaddb <= "111010010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101010";
				elsif cntr ="000111101010" THEN
				      ioadda <= "011010101";
				      ioaddb <= "111010100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101011";
				elsif cntr ="000111101011" THEN
				      ioadda <= "011010111";
				      ioaddb <= "111010110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101100";
				elsif cntr ="000111101100" THEN
				      ioadda <= "011011001";
				      ioaddb <= "111011000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101101";
				elsif cntr ="000111101101" THEN
				      ioadda <= "011011011";
				      ioaddb <= "111011010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101110";
				elsif cntr ="000111101110" THEN
				      ioadda <= "011011101";
				      ioaddb <= "111011100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111101111";
				elsif cntr ="000111101111" THEN
				      ioadda <= "011011111";
				      ioaddb <= "111011110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110000";
				elsif cntr ="000111110000" THEN
				      ioadda <= "011100001";
				      ioaddb <= "111100000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110001";
				elsif cntr ="000111110001" THEN
				      ioadda <= "011100011";
				      ioaddb <= "111100010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110010";
				elsif cntr ="000111110010" THEN
				      ioadda <= "011100101";
				      ioaddb <= "111100100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110011";
				elsif cntr ="000111110011" THEN
				      ioadda <= "011100111";
				      ioaddb <= "111100110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110100";
				elsif cntr ="000111110100" THEN
				      ioadda <= "011101001";
				      ioaddb <= "111101000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110101";
				elsif cntr ="000111110101" THEN
				      ioadda <= "011101011";
				      ioaddb <= "111101010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110110";
				elsif cntr ="000111110110" THEN
				      ioadda <= "011101101";
				      ioaddb <= "111101100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111110111";
				elsif cntr ="000111110111" THEN
				      ioadda <= "011101111";
				      ioaddb <= "111101110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111000";
				elsif cntr ="000111111000" THEN
				      ioadda <= "011110001";
				      ioaddb <= "111110000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111001";
				elsif cntr ="000111111001" THEN
				      ioadda <= "011110011";
				      ioaddb <= "111110010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111010";
				elsif cntr ="000111111010" THEN
				      ioadda <= "011110101";
				      ioaddb <= "111110100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111011";
				elsif cntr ="000111111011" THEN
				      ioadda <= "011110111";
				      ioaddb <= "111110110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111100";
				elsif cntr ="000111111100" THEN
				      ioadda <= "011111001";
				      ioaddb <= "111111000";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111101";
				elsif cntr ="000111111101" THEN
				      ioadda <= "011111011";
				      ioaddb <= "111111010";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111110";
				elsif cntr ="000111111110" THEN
				      ioadda <= "011111101";
				      ioaddb <= "111111100";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "000111111111";
				elsif cntr ="000111111111" THEN
				      ioadda <= "011111111";
				      ioaddb <= "111111110";
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000000000";
				elsif cntr ="001000000000" THEN	
				      t1addb <= "00000000";      
				      zetain <= "01000000";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000000001";
				elsif cntr ="001000000001" THEN	
				      t1addb <= "00000001";      
				      zetain <= "11000000";      
				      bfrjin   <= iodouta;
				      bfrjplin <= iodoutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000000010";
				elsif cntr ="001000000010" THEN	
				      t1addb <= "00000010";      
				      zetain <= "01000001";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				            
				            
				            
				      cntr <= "001000000011";      
				elsif cntr ="001000000011" THEN	      
				      t1addb <= "00000011";      
				      zetain <= "11000001";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001000000100";            
				elsif cntr ="001000000100" THEN	         
				      t1addb <= "00000100";      
				      zetain <= "01000010";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001000000101";               
				elsif cntr ="001000000101" THEN	            
				      t1addb <= "00000101";      
				      zetain <= "11000010";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001000000110";            
				elsif cntr ="001000000110" THEN	         
				      t1addb <= "00000110";      
				      zetain <= "01000011";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001000000111";                  
				elsif cntr ="001000000111" THEN	               
				      t1addb <= "00000111";      
				      zetain <= "11000011";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= zetaout;      
				      
				      
				      
				                                  
				                                  
				                                  
				      cntr <= "001000001000";     
				elsif cntr ="001000001000" THEN	  
				      t1addb <= "00001000";
				      zetain <= "01000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				
				
				
				      
				      
				      
				      cntr <= "001000001001";
				elsif cntr ="001000001001" THEN
				      t1addb <= "00001001";
				      zetain <= "11000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001010";
				elsif cntr ="001000001010" THEN
				      t1addb <= "00001010";
				      zetain <= "01000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001011";
				elsif cntr ="001000001011" THEN
				      t1addb <= "00001011";
				      zetain <= "11000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001100";
				elsif cntr ="001000001100" THEN
				      t1addb <= "00001100";
				      zetain <= "01000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001101";
				elsif cntr ="001000001101" THEN
				      t1addb <= "00001101";
				      zetain <= "11000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001110";
				elsif cntr ="001000001110" THEN
				      t1addb <= "00001110";
				      zetain <= "01000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000001111";
				elsif cntr ="001000001111" THEN
				      t1addb <= "00001111";
				      zetain <= "11000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010000";
				elsif cntr ="001000010000" THEN
				      t1addb <= "00010000";
				      zetain <= "01001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010001";
				elsif cntr ="001000010001" THEN
				      t1addb <= "00010001";
				      zetain <= "11001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010010";
				elsif cntr ="001000010010" THEN
				      t1addb <= "00010010";
				      zetain <= "01001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010011";
				elsif cntr ="001000010011" THEN
				      t1addb <= "00010011";
				      zetain <= "11001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010100";
				elsif cntr ="001000010100" THEN
				      t1addb <= "00010100";
				      zetain <= "01001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010101";
				elsif cntr ="001000010101" THEN
				      t1addb <= "00010101";
				      zetain <= "11001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010110";
				elsif cntr ="001000010110" THEN
				      t1addb <= "00010110";
				      zetain <= "01001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000010111";
				elsif cntr ="001000010111" THEN
				      t1addb <= "00010111";
				      zetain <= "11001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011000";
				elsif cntr ="001000011000" THEN
				      t1addb <= "00011000";
				      zetain <= "01001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011001";
				elsif cntr ="001000011001" THEN
				      t1addb <= "00011001";
				      zetain <= "11001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011010";
				elsif cntr ="001000011010" THEN
				      t1addb <= "00011010";
				      zetain <= "01001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011011";
				elsif cntr ="001000011011" THEN
				      t1addb <= "00011011";
				      zetain <= "11001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011100";
				elsif cntr ="001000011100" THEN
				      t1addb <= "00011100";
				      zetain <= "01001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011101";
				elsif cntr ="001000011101" THEN
				      t1addb <= "00011101";
				      zetain <= "11001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011110";
				elsif cntr ="001000011110" THEN
				      t1addb <= "00011110";
				      zetain <= "01001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000011111";
				elsif cntr ="001000011111" THEN
				      t1addb <= "00011111";
				      zetain <= "11001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100000";
				elsif cntr ="001000100000" THEN
				      t1addb <= "00100000";
				      zetain <= "01010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100001";
				elsif cntr ="001000100001" THEN
				      t1addb <= "00100001";
				      zetain <= "11010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100010";
				elsif cntr ="001000100010" THEN
				      t1addb <= "00100010";
				      zetain <= "01010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100011";
				elsif cntr ="001000100011" THEN
				      t1addb <= "00100011";
				      zetain <= "11010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100100";
				elsif cntr ="001000100100" THEN
				      t1addb <= "00100100";
				      zetain <= "01010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100101";
				elsif cntr ="001000100101" THEN
				      t1addb <= "00100101";
				      zetain <= "11010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100110";
				elsif cntr ="001000100110" THEN
				      t1addb <= "00100110";
				      zetain <= "01010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000100111";
				elsif cntr ="001000100111" THEN
				      t1addb <= "00100111";
				      zetain <= "11010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101000";
				elsif cntr ="001000101000" THEN
				      t1addb <= "00101000";
				      zetain <= "01010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101001";
				elsif cntr ="001000101001" THEN
				      t1addb <= "00101001";
				      zetain <= "11010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101010";
				elsif cntr ="001000101010" THEN
				      t1addb <= "00101010";
				      zetain <= "01010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101011";
				elsif cntr ="001000101011" THEN
				      t1addb <= "00101011";
				      zetain <= "11010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101100";
				elsif cntr ="001000101100" THEN
				      t1addb <= "00101100";
				      zetain <= "01010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101101";
				elsif cntr ="001000101101" THEN
				      t1addb <= "00101101";
				      zetain <= "11010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101110";
				elsif cntr ="001000101110" THEN
				      t1addb <= "00101110";
				      zetain <= "01010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000101111";
				elsif cntr ="001000101111" THEN
				      t1addb <= "00101111";
				      zetain <= "11010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110000";
				elsif cntr ="001000110000" THEN
				      t1addb <= "00110000";
				      zetain <= "01011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110001";
				elsif cntr ="001000110001" THEN
				      t1addb <= "00110001";
				      zetain <= "11011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110010";
				elsif cntr ="001000110010" THEN
				      t1addb <= "00110010";
				      zetain <= "01011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110011";
				elsif cntr ="001000110011" THEN
				      t1addb <= "00110011";
				      zetain <= "11011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110100";
				elsif cntr ="001000110100" THEN
				      t1addb <= "00110100";
				      zetain <= "01011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110101";
				elsif cntr ="001000110101" THEN
				      t1addb <= "00110101";
				      zetain <= "11011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110110";
				elsif cntr ="001000110110" THEN
				      t1addb <= "00110110";
				      zetain <= "01011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000110111";
				elsif cntr ="001000110111" THEN
				      t1addb <= "00110111";
				      zetain <= "11011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111000";
				elsif cntr ="001000111000" THEN
				      t1addb <= "00111000";
				      zetain <= "01011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111001";
				elsif cntr ="001000111001" THEN
				      t1addb <= "00111001";
				      zetain <= "11011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111010";
				elsif cntr ="001000111010" THEN
				      t1addb <= "00111010";
				      zetain <= "01011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111011";
				elsif cntr ="001000111011" THEN
				      t1addb <= "00111011";
				      zetain <= "11011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111100";
				elsif cntr ="001000111100" THEN
				      t1addb <= "00111100";
				      zetain <= "01011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111101";
				elsif cntr ="001000111101" THEN
				      t1addb <= "00111101";
				      zetain <= "11011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111110";
				elsif cntr ="001000111110" THEN
				      t1addb <= "00111110";
				      zetain <= "01011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001000111111";
				elsif cntr ="001000111111" THEN
				      t1addb <= "00111111";
				      zetain <= "11011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000000";
				elsif cntr ="001001000000" THEN
				      t1addb <= "01000000";
				      zetain <= "01100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000001";
				elsif cntr ="001001000001" THEN
				      t1addb <= "01000001";
				      zetain <= "11100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000010";
				elsif cntr ="001001000010" THEN
				      t1addb <= "01000010";
				      zetain <= "01100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000011";
				elsif cntr ="001001000011" THEN
				      t1addb <= "01000011";
				      zetain <= "11100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000100";
				elsif cntr ="001001000100" THEN
				      t1addb <= "01000100";
				      zetain <= "01100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000101";
				elsif cntr ="001001000101" THEN
				      t1addb <= "01000101";
				      zetain <= "11100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000110";
				elsif cntr ="001001000110" THEN
				      t1addb <= "01000110";
				      zetain <= "01100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001000111";
				elsif cntr ="001001000111" THEN
				      t1addb <= "01000111";
				      zetain <= "11100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001000";
				elsif cntr ="001001001000" THEN
				      t1addb <= "01001000";
				      zetain <= "01100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001001";
				elsif cntr ="001001001001" THEN
				      t1addb <= "01001001";
				      zetain <= "11100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001010";
				elsif cntr ="001001001010" THEN
				      t1addb <= "01001010";
				      zetain <= "01100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001011";
				elsif cntr ="001001001011" THEN
				      t1addb <= "01001011";
				      zetain <= "11100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001100";
				elsif cntr ="001001001100" THEN
				      t1addb <= "01001100";
				      zetain <= "01100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001101";
				elsif cntr ="001001001101" THEN
				      t1addb <= "01001101";
				      zetain <= "11100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001110";
				elsif cntr ="001001001110" THEN
				      t1addb <= "01001110";
				      zetain <= "01100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001001111";
				elsif cntr ="001001001111" THEN
				      t1addb <= "01001111";
				      zetain <= "11100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010000";
				elsif cntr ="001001010000" THEN
				      t1addb <= "01010000";
				      zetain <= "01101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010001";
				elsif cntr ="001001010001" THEN
				      t1addb <= "01010001";
				      zetain <= "11101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010010";
				elsif cntr ="001001010010" THEN
				      t1addb <= "01010010";
				      zetain <= "01101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010011";
				elsif cntr ="001001010011" THEN
				      t1addb <= "01010011";
				      zetain <= "11101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010100";
				elsif cntr ="001001010100" THEN
				      t1addb <= "01010100";
				      zetain <= "01101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010101";
				elsif cntr ="001001010101" THEN
				      t1addb <= "01010101";
				      zetain <= "11101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010110";
				elsif cntr ="001001010110" THEN
				      t1addb <= "01010110";
				      zetain <= "01101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001010111";
				elsif cntr ="001001010111" THEN
				      t1addb <= "01010111";
				      zetain <= "11101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011000";
				elsif cntr ="001001011000" THEN
				      t1addb <= "01011000";
				      zetain <= "01101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011001";
				elsif cntr ="001001011001" THEN
				      t1addb <= "01011001";
				      zetain <= "11101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011010";
				elsif cntr ="001001011010" THEN
				      t1addb <= "01011010";
				      zetain <= "01101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011011";
				elsif cntr ="001001011011" THEN
				      t1addb <= "01011011";
				      zetain <= "11101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011100";
				elsif cntr ="001001011100" THEN
				      t1addb <= "01011100";
				      zetain <= "01101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011101";
				elsif cntr ="001001011101" THEN
				      t1addb <= "01011101";
				      zetain <= "11101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011110";
				elsif cntr ="001001011110" THEN
				      t1addb <= "01011110";
				      zetain <= "01101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001011111";
				elsif cntr ="001001011111" THEN
				      t1addb <= "01011111";
				      zetain <= "11101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100000";
				elsif cntr ="001001100000" THEN
				      t1addb <= "01100000";
				      zetain <= "01110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100001";
				elsif cntr ="001001100001" THEN
				      t1addb <= "01100001";
				      zetain <= "11110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100010";
				elsif cntr ="001001100010" THEN
				      t1addb <= "01100010";
				      zetain <= "01110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100011";
				elsif cntr ="001001100011" THEN
				      t1addb <= "01100011";
				      zetain <= "11110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100100";
				elsif cntr ="001001100100" THEN
				      t1addb <= "01100100";
				      zetain <= "01110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100101";
				elsif cntr ="001001100101" THEN
				      t1addb <= "01100101";
				      zetain <= "11110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100110";
				elsif cntr ="001001100110" THEN
				      t1addb <= "01100110";
				      zetain <= "01110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001100111";
				elsif cntr ="001001100111" THEN
				      t1addb <= "01100111";
				      zetain <= "11110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101000";
				elsif cntr ="001001101000" THEN
				      t1addb <= "01101000";
				      zetain <= "01110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101001";
				elsif cntr ="001001101001" THEN
				      t1addb <= "01101001";
				      zetain <= "11110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101010";
				elsif cntr ="001001101010" THEN
				      t1addb <= "01101010";
				      zetain <= "01110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101011";
				elsif cntr ="001001101011" THEN
				      t1addb <= "01101011";
				      zetain <= "11110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101100";
				elsif cntr ="001001101100" THEN
				      t1addb <= "01101100";
				      zetain <= "01110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101101";
				elsif cntr ="001001101101" THEN
				      t1addb <= "01101101";
				      zetain <= "11110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101110";
				elsif cntr ="001001101110" THEN
				      t1addb <= "01101110";
				      zetain <= "01110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001101111";
				elsif cntr ="001001101111" THEN
				      t1addb <= "01101111";
				      zetain <= "11110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110000";
				elsif cntr ="001001110000" THEN
				      t1addb <= "01110000";
				      zetain <= "01111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110001";
				elsif cntr ="001001110001" THEN
				      t1addb <= "01110001";
				      zetain <= "11111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110010";
				elsif cntr ="001001110010" THEN
				      t1addb <= "01110010";
				      zetain <= "01111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110011";
				elsif cntr ="001001110011" THEN
				      t1addb <= "01110011";
				      zetain <= "11111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110100";
				elsif cntr ="001001110100" THEN
				      t1addb <= "01110100";
				      zetain <= "01111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110101";
				elsif cntr ="001001110101" THEN
				      t1addb <= "01110101";
				      zetain <= "11111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110110";
				elsif cntr ="001001110110" THEN
				      t1addb <= "01110110";
				      zetain <= "01111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001110111";
				elsif cntr ="001001110111" THEN
				      t1addb <= "01110111";
				      zetain <= "11111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111000";
				elsif cntr ="001001111000" THEN
				      t1addb <= "01111000";
				      zetain <= "01111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111001";
				elsif cntr ="001001111001" THEN
				      t1addb <= "01111001";
				      zetain <= "11111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111010";
				elsif cntr ="001001111010" THEN
				      t1addb <= "01111010";
				      zetain <= "01111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111011";
				elsif cntr ="001001111011" THEN
				      t1addb <= "01111011";
				      zetain <= "11111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111100";
				elsif cntr ="001001111100" THEN
				      t1addb <= "01111100";
				      zetain <= "01111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111101";
				elsif cntr ="001001111101" THEN
				      t1addb <= "01111101";
				      zetain <= "11111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111110";
				elsif cntr ="001001111110" THEN
				      t1addb <= "01111110";
				      zetain <= "01111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001001111111";
				elsif cntr ="001001111111" THEN
				      t1addb <= "01111111";
				      zetain <= "11111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010000000";
				elsif cntr ="001010000000" THEN
				      
				      
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010000001";
				elsif cntr ="001010000001" THEN
				      
				      
				      bfrjin   <= t1doutb;
				      bfrjplin <= zetaout;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010000010";
				elsif cntr ="001010000010" THEN
				      
				      
				      
				      
				      
				      
				      
				            
				            
				            
				      cntr <= "001010000011";      
				elsif cntr ="001010000011" THEN      
				      
				      
				      
				      
				      
				      
				      
				                  
				                  
				                  
				      cntr <= "001010000100";            
				elsif cntr ="001010000100" THEN            
				      
				      
				      
				      
				      
				      
				      
				                        
				                        
				                        
				      cntr <= "001010000101";             
				elsif cntr ="001010000101" THEN           
				      
				      
				      
				      
				      
				      
				      
				                              
				                              
				                              
				      cntr <= "001010000110";         
				elsif cntr ="001010000110" THEN       
				      
				      
				      
				      
				      
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001010000111";             
				elsif cntr ="001010000111" THEN           
				      t1addb <= "00000000";      
				      t2addb <= "00000000";      
				      
				      
				    
				      
				      
				                                    
				                                    
				                                    
				      cntr <= "001010001000";         
				elsif cntr ="001010001000" THEN       
				      t1addb <= "00000001";
				      t2addb <= "00000001";
				
				
				
				 	 bfmod <="11";
				
				
				
				
				
				
				
				
				
				
				      cntr <= "001010001001";
				elsif cntr ="001010001001" THEN
				      t1addb <= "00000010";
				      t2addb <= "00000010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				
				
				
				
				
				
				
				
				
				      cntr <= "001010001010";
				elsif cntr ="001010001010" THEN
				      t1addb <= "00000011";
				      t2addb <= "00000011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "001010001011";
				elsif cntr ="001010001011" THEN
				      t1addb <= "00000100";
				      t2addb <= "00000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001100";
				elsif cntr ="001010001100" THEN
				      t1addb <= "00000101";
				      t2addb <= "00000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001101";
				elsif cntr ="001010001101" THEN
				      t1addb <= "00000110";
				      t2addb <= "00000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001110";
				elsif cntr ="001010001110" THEN
				      t1addb <= "00000111";
				      t2addb <= "00000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010001111";
				elsif cntr ="001010001111" THEN
				      t1addb <= "00001000";
				      t2addb <= "00001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010000";
				elsif cntr ="001010010000" THEN
				      t1addb <= "00001001";
				      t2addb <= "00001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010001";
				elsif cntr ="001010010001" THEN
				      t1addb <= "00001010";
				      t2addb <= "00001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010010";
				elsif cntr ="001010010010" THEN
				      t1addb <= "00001011";
				      t2addb <= "00001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010011";
				elsif cntr ="001010010011" THEN
				      t1addb <= "00001100";
				      t2addb <= "00001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010100";
				elsif cntr ="001010010100" THEN
				      t1addb <= "00001101";
				      t2addb <= "00001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010101";
				elsif cntr ="001010010101" THEN
				      t1addb <= "00001110";
				      t2addb <= "00001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010110";
				elsif cntr ="001010010110" THEN
				      t1addb <= "00001111";
				      t2addb <= "00001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010010111";
				elsif cntr ="001010010111" THEN
				      t1addb <= "00010000";
				      t2addb <= "00010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011000";
				elsif cntr ="001010011000" THEN
				      t1addb <= "00010001";
				      t2addb <= "00010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011001";
				elsif cntr ="001010011001" THEN
				      t1addb <= "00010010";
				      t2addb <= "00010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011010";
				elsif cntr ="001010011010" THEN
				      t1addb <= "00010011";
				      t2addb <= "00010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011011";
				elsif cntr ="001010011011" THEN
				      t1addb <= "00010100";
				      t2addb <= "00010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011100";
				elsif cntr ="001010011100" THEN
				      t1addb <= "00010101";
				      t2addb <= "00010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011101";
				elsif cntr ="001010011101" THEN
				      t1addb <= "00010110";
				      t2addb <= "00010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011110";
				elsif cntr ="001010011110" THEN
				      t1addb <= "00010111";
				      t2addb <= "00010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010011111";
				elsif cntr ="001010011111" THEN
				      t1addb <= "00011000";
				      t2addb <= "00011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100000";
				elsif cntr ="001010100000" THEN
				      t1addb <= "00011001";
				      t2addb <= "00011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100001";
				elsif cntr ="001010100001" THEN
				      t1addb <= "00011010";
				      t2addb <= "00011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100010";
				elsif cntr ="001010100010" THEN
				      t1addb <= "00011011";
				      t2addb <= "00011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100011";
				elsif cntr ="001010100011" THEN
				      t1addb <= "00011100";
				      t2addb <= "00011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100100";
				elsif cntr ="001010100100" THEN
				      t1addb <= "00011101";
				      t2addb <= "00011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100101";
				elsif cntr ="001010100101" THEN
				      t1addb <= "00011110";
				      t2addb <= "00011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100110";
				elsif cntr ="001010100110" THEN
				      t1addb <= "00011111";
				      t2addb <= "00011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010100111";
				elsif cntr ="001010100111" THEN
				      t1addb <= "00100000";
				      t2addb <= "00100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101000";
				elsif cntr ="001010101000" THEN
				      t1addb <= "00100001";
				      t2addb <= "00100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101001";
				elsif cntr ="001010101001" THEN
				      t1addb <= "00100010";
				      t2addb <= "00100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101010";
				elsif cntr ="001010101010" THEN
				      t1addb <= "00100011";
				      t2addb <= "00100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101011";
				elsif cntr ="001010101011" THEN
				      t1addb <= "00100100";
				      t2addb <= "00100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101100";
				elsif cntr ="001010101100" THEN
				      t1addb <= "00100101";
				      t2addb <= "00100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101101";
				elsif cntr ="001010101101" THEN
				      t1addb <= "00100110";
				      t2addb <= "00100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101110";
				elsif cntr ="001010101110" THEN
				      t1addb <= "00100111";
				      t2addb <= "00100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010101111";
				elsif cntr ="001010101111" THEN
				      t1addb <= "00101000";
				      t2addb <= "00101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110000";
				elsif cntr ="001010110000" THEN
				      t1addb <= "00101001";
				      t2addb <= "00101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110001";
				elsif cntr ="001010110001" THEN
				      t1addb <= "00101010";
				      t2addb <= "00101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110010";
				elsif cntr ="001010110010" THEN
				      t1addb <= "00101011";
				      t2addb <= "00101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110011";
				elsif cntr ="001010110011" THEN
				      t1addb <= "00101100";
				      t2addb <= "00101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110100";
				elsif cntr ="001010110100" THEN
				      t1addb <= "00101101";
				      t2addb <= "00101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110101";
				elsif cntr ="001010110101" THEN
				      t1addb <= "00101110";
				      t2addb <= "00101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110110";
				elsif cntr ="001010110110" THEN
				      t1addb <= "00101111";
				      t2addb <= "00101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010110111";
				elsif cntr ="001010110111" THEN
				      t1addb <= "00110000";
				      t2addb <= "00110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111000";
				elsif cntr ="001010111000" THEN
				      t1addb <= "00110001";
				      t2addb <= "00110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111001";
				elsif cntr ="001010111001" THEN
				      t1addb <= "00110010";
				      t2addb <= "00110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111010";
				elsif cntr ="001010111010" THEN
				      t1addb <= "00110011";
				      t2addb <= "00110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111011";
				elsif cntr ="001010111011" THEN
				      t1addb <= "00110100";
				      t2addb <= "00110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111100";
				elsif cntr ="001010111100" THEN
				      t1addb <= "00110101";
				      t2addb <= "00110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111101";
				elsif cntr ="001010111101" THEN
				      t1addb <= "00110110";
				      t2addb <= "00110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111110";
				elsif cntr ="001010111110" THEN
				      t1addb <= "00110111";
				      t2addb <= "00110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001010111111";
				elsif cntr ="001010111111" THEN
				      t1addb <= "00111000";
				      t2addb <= "00111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000000";
				elsif cntr ="001011000000" THEN
				      t1addb <= "00111001";
				      t2addb <= "00111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000001";
				elsif cntr ="001011000001" THEN
				      t1addb <= "00111010";
				      t2addb <= "00111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000010";
				elsif cntr ="001011000010" THEN
				      t1addb <= "00111011";
				      t2addb <= "00111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000011";
				elsif cntr ="001011000011" THEN
				      t1addb <= "00111100";
				      t2addb <= "00111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000100";
				elsif cntr ="001011000100" THEN
				      t1addb <= "00111101";
				      t2addb <= "00111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000101";
				elsif cntr ="001011000101" THEN
				      t1addb <= "00111110";
				      t2addb <= "00111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000110";
				elsif cntr ="001011000110" THEN
				      t1addb <= "00111111";
				      t2addb <= "00111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011000111";
				elsif cntr ="001011000111" THEN
				      t1addb <= "01000000";
				      t2addb <= "01000000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001000";
				elsif cntr ="001011001000" THEN
				      t1addb <= "01000001";
				      t2addb <= "01000001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001001";
				elsif cntr ="001011001001" THEN
				      t1addb <= "01000010";
				      t2addb <= "01000010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001010";
				elsif cntr ="001011001010" THEN
				      t1addb <= "01000011";
				      t2addb <= "01000011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001011";
				elsif cntr ="001011001011" THEN
				      t1addb <= "01000100";
				      t2addb <= "01000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001100";
				elsif cntr ="001011001100" THEN
				      t1addb <= "01000101";
				      t2addb <= "01000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001101";
				elsif cntr ="001011001101" THEN
				      t1addb <= "01000110";
				      t2addb <= "01000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001110";
				elsif cntr ="001011001110" THEN
				      t1addb <= "01000111";
				      t2addb <= "01000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011001111";
				elsif cntr ="001011001111" THEN
				      t1addb <= "01001000";
				      t2addb <= "01001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010000";
				elsif cntr ="001011010000" THEN
				      t1addb <= "01001001";
				      t2addb <= "01001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010001";
				elsif cntr ="001011010001" THEN
				      t1addb <= "01001010";
				      t2addb <= "01001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010010";
				elsif cntr ="001011010010" THEN
				      t1addb <= "01001011";
				      t2addb <= "01001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010011";
				elsif cntr ="001011010011" THEN
				      t1addb <= "01001100";
				      t2addb <= "01001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010100";
				elsif cntr ="001011010100" THEN
				      t1addb <= "01001101";
				      t2addb <= "01001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010101";
				elsif cntr ="001011010101" THEN
				      t1addb <= "01001110";
				      t2addb <= "01001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010110";
				elsif cntr ="001011010110" THEN
				      t1addb <= "01001111";
				      t2addb <= "01001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011010111";
				elsif cntr ="001011010111" THEN
				      t1addb <= "01010000";
				      t2addb <= "01010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011000";
				elsif cntr ="001011011000" THEN
				      t1addb <= "01010001";
				      t2addb <= "01010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011001";
				elsif cntr ="001011011001" THEN
				      t1addb <= "01010010";
				      t2addb <= "01010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011010";
				elsif cntr ="001011011010" THEN
				      t1addb <= "01010011";
				      t2addb <= "01010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011011";
				elsif cntr ="001011011011" THEN
				      t1addb <= "01010100";
				      t2addb <= "01010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011100";
				elsif cntr ="001011011100" THEN
				      t1addb <= "01010101";
				      t2addb <= "01010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011101";
				elsif cntr ="001011011101" THEN
				      t1addb <= "01010110";
				      t2addb <= "01010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011110";
				elsif cntr ="001011011110" THEN
				      t1addb <= "01010111";
				      t2addb <= "01010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011011111";
				elsif cntr ="001011011111" THEN
				      t1addb <= "01011000";
				      t2addb <= "01011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100000";
				elsif cntr ="001011100000" THEN
				      t1addb <= "01011001";
				      t2addb <= "01011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100001";
				elsif cntr ="001011100001" THEN
				      t1addb <= "01011010";
				      t2addb <= "01011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100010";
				elsif cntr ="001011100010" THEN
				      t1addb <= "01011011";
				      t2addb <= "01011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100011";
				elsif cntr ="001011100011" THEN
				      t1addb <= "01011100";
				      t2addb <= "01011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100100";
				elsif cntr ="001011100100" THEN
				      t1addb <= "01011101";
				      t2addb <= "01011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100101";
				elsif cntr ="001011100101" THEN
				      t1addb <= "01011110";
				      t2addb <= "01011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100110";
				elsif cntr ="001011100110" THEN
				      t1addb <= "01011111";
				      t2addb <= "01011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011100111";
				elsif cntr ="001011100111" THEN
				      t1addb <= "01100000";
				      t2addb <= "01100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101000";
				elsif cntr ="001011101000" THEN
				      t1addb <= "01100001";
				      t2addb <= "01100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101001";
				elsif cntr ="001011101001" THEN
				      t1addb <= "01100010";
				      t2addb <= "01100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101010";
				elsif cntr ="001011101010" THEN
				      t1addb <= "01100011";
				      t2addb <= "01100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101011";
				elsif cntr ="001011101011" THEN
				      t1addb <= "01100100";
				      t2addb <= "01100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101100";
				elsif cntr ="001011101100" THEN
				      t1addb <= "01100101";
				      t2addb <= "01100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101101";
				elsif cntr ="001011101101" THEN
				      t1addb <= "01100110";
				      t2addb <= "01100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101110";
				elsif cntr ="001011101110" THEN
				      t1addb <= "01100111";
				      t2addb <= "01100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011101111";
				elsif cntr ="001011101111" THEN
				      t1addb <= "01101000";
				      t2addb <= "01101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110000";
				elsif cntr ="001011110000" THEN
				      t1addb <= "01101001";
				      t2addb <= "01101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110001";
				elsif cntr ="001011110001" THEN
				      t1addb <= "01101010";
				      t2addb <= "01101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110010";
				elsif cntr ="001011110010" THEN
				      t1addb <= "01101011";
				      t2addb <= "01101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110011";
				elsif cntr ="001011110011" THEN
				      t1addb <= "01101100";
				      t2addb <= "01101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110100";
				elsif cntr ="001011110100" THEN
				      t1addb <= "01101101";
				      t2addb <= "01101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110101";
				elsif cntr ="001011110101" THEN
				      t1addb <= "01101110";
				      t2addb <= "01101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110110";
				elsif cntr ="001011110110" THEN
				      t1addb <= "01101111";
				      t2addb <= "01101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011110111";
				elsif cntr ="001011110111" THEN
				      t1addb <= "01110000";
				      t2addb <= "01110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111000";
				elsif cntr ="001011111000" THEN
				      t1addb <= "01110001";
				      t2addb <= "01110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111001";
				elsif cntr ="001011111001" THEN
				      t1addb <= "01110010";
				      t2addb <= "01110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111010";
				elsif cntr ="001011111010" THEN
				      t1addb <= "01110011";
				      t2addb <= "01110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111011";
				elsif cntr ="001011111011" THEN
				      t1addb <= "01110100";
				      t2addb <= "01110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111100";
				elsif cntr ="001011111100" THEN
				      t1addb <= "01110101";
				      t2addb <= "01110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111101";
				elsif cntr ="001011111101" THEN
				      t1addb <= "01110110";
				      t2addb <= "01110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111110";
				elsif cntr ="001011111110" THEN
				      t1addb <= "01110111";
				      t2addb <= "01110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001011111111";
				elsif cntr ="001011111111" THEN
				      t1addb <= "01111000";
				      t2addb <= "01111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000000";
				elsif cntr ="001100000000" THEN
				      t1addb <= "01111001";
				      t2addb <= "01111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000001";
				elsif cntr ="001100000001" THEN
				      t1addb <= "01111010";
				      t2addb <= "01111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000010";
				elsif cntr ="001100000010" THEN
				      t1addb <= "01111011";
				      t2addb <= "01111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000011";
				elsif cntr ="001100000011" THEN
				      t1addb <= "01111100";
				      t2addb <= "01111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000100";
				elsif cntr ="001100000100" THEN
				      t1addb <= "01111101";
				      t2addb <= "01111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000101";
				elsif cntr ="001100000101" THEN
				      t1addb <= "01111110";
				      t2addb <= "01111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000110";
				elsif cntr ="001100000110" THEN
				      t1addb <= "01111111";
				      t2addb <= "01111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100000111";
				elsif cntr ="001100000111" THEN
				      t1addb <= "10000000";      
				      t2addb <= "10000000";      
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001000";
				elsif cntr ="001100001000" THEN
				      t1addb <= "10000001";      
				      t2addb <= "10000001";      
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001001";
				elsif cntr ="001100001001" THEN
				      t1addb <= "10000010";      
				      t2addb <= "10000010";      
				      bfrjin   <= t1doutb;      
				      bfrjplin <= t2doutb;      
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001010";
				elsif cntr ="001100001010" THEN
				      t1addb <= "10000011";
				      t2addb <= "10000011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				
				
				
				      
				      
				      
				      cntr <= "001100001011";
				elsif cntr ="001100001011" THEN
				      t1addb <= "10000100";
				      t2addb <= "10000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001100";
				elsif cntr ="001100001100" THEN
				      t1addb <= "10000101";
				      t2addb <= "10000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001101";
				elsif cntr ="001100001101" THEN
				      t1addb <= "10000110";
				      t2addb <= "10000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001110";
				elsif cntr ="001100001110" THEN
				      t1addb <= "10000111";
				      t2addb <= "10000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100001111";
				elsif cntr ="001100001111" THEN
				      t1addb <= "10001000";
				      t2addb <= "10001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010000";
				elsif cntr ="001100010000" THEN
				      t1addb <= "10001001";
				      t2addb <= "10001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010001";
				elsif cntr ="001100010001" THEN
				      t1addb <= "10001010";
				      t2addb <= "10001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010010";
				elsif cntr ="001100010010" THEN
				      t1addb <= "10001011";
				      t2addb <= "10001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010011";
				elsif cntr ="001100010011" THEN
				      t1addb <= "10001100";
				      t2addb <= "10001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010100";
				elsif cntr ="001100010100" THEN
				      t1addb <= "10001101";
				      t2addb <= "10001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010101";
				elsif cntr ="001100010101" THEN
				      t1addb <= "10001110";
				      t2addb <= "10001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010110";
				elsif cntr ="001100010110" THEN
				      t1addb <= "10001111";
				      t2addb <= "10001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100010111";
				elsif cntr ="001100010111" THEN
				      t1addb <= "10010000";
				      t2addb <= "10010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011000";
				elsif cntr ="001100011000" THEN
				      t1addb <= "10010001";
				      t2addb <= "10010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011001";
				elsif cntr ="001100011001" THEN
				      t1addb <= "10010010";
				      t2addb <= "10010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011010";
				elsif cntr ="001100011010" THEN
				      t1addb <= "10010011";
				      t2addb <= "10010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011011";
				elsif cntr ="001100011011" THEN
				      t1addb <= "10010100";
				      t2addb <= "10010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011100";
				elsif cntr ="001100011100" THEN
				      t1addb <= "10010101";
				      t2addb <= "10010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011101";
				elsif cntr ="001100011101" THEN
				      t1addb <= "10010110";
				      t2addb <= "10010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011110";
				elsif cntr ="001100011110" THEN
				      t1addb <= "10010111";
				      t2addb <= "10010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100011111";
				elsif cntr ="001100011111" THEN
				      t1addb <= "10011000";
				      t2addb <= "10011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100000";
				elsif cntr ="001100100000" THEN
				      t1addb <= "10011001";
				      t2addb <= "10011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100001";
				elsif cntr ="001100100001" THEN
				      t1addb <= "10011010";
				      t2addb <= "10011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100010";
				elsif cntr ="001100100010" THEN
				      t1addb <= "10011011";
				      t2addb <= "10011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100011";
				elsif cntr ="001100100011" THEN
				      t1addb <= "10011100";
				      t2addb <= "10011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100100";
				elsif cntr ="001100100100" THEN
				      t1addb <= "10011101";
				      t2addb <= "10011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100101";
				elsif cntr ="001100100101" THEN
				      t1addb <= "10011110";
				      t2addb <= "10011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100110";
				elsif cntr ="001100100110" THEN
				      t1addb <= "10011111";
				      t2addb <= "10011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100100111";
				elsif cntr ="001100100111" THEN
				      t1addb <= "10100000";
				      t2addb <= "10100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101000";
				elsif cntr ="001100101000" THEN
				      t1addb <= "10100001";
				      t2addb <= "10100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101001";
				elsif cntr ="001100101001" THEN
				      t1addb <= "10100010";
				      t2addb <= "10100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101010";
				elsif cntr ="001100101010" THEN
				      t1addb <= "10100011";
				      t2addb <= "10100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101011";
				elsif cntr ="001100101011" THEN
				      t1addb <= "10100100";
				      t2addb <= "10100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101100";
				elsif cntr ="001100101100" THEN
				      t1addb <= "10100101";
				      t2addb <= "10100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101101";
				elsif cntr ="001100101101" THEN
				      t1addb <= "10100110";
				      t2addb <= "10100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101110";
				elsif cntr ="001100101110" THEN
				      t1addb <= "10100111";
				      t2addb <= "10100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100101111";
				elsif cntr ="001100101111" THEN
				      t1addb <= "10101000";
				      t2addb <= "10101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110000";
				elsif cntr ="001100110000" THEN
				      t1addb <= "10101001";
				      t2addb <= "10101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110001";
				elsif cntr ="001100110001" THEN
				      t1addb <= "10101010";
				      t2addb <= "10101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110010";
				elsif cntr ="001100110010" THEN
				      t1addb <= "10101011";
				      t2addb <= "10101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110011";
				elsif cntr ="001100110011" THEN
				      t1addb <= "10101100";
				      t2addb <= "10101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110100";
				elsif cntr ="001100110100" THEN
				      t1addb <= "10101101";
				      t2addb <= "10101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110101";
				elsif cntr ="001100110101" THEN
				      t1addb <= "10101110";
				      t2addb <= "10101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110110";
				elsif cntr ="001100110110" THEN
				      t1addb <= "10101111";
				      t2addb <= "10101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100110111";
				elsif cntr ="001100110111" THEN
				      t1addb <= "10110000";
				      t2addb <= "10110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111000";
				elsif cntr ="001100111000" THEN
				      t1addb <= "10110001";
				      t2addb <= "10110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111001";
				elsif cntr ="001100111001" THEN
				      t1addb <= "10110010";
				      t2addb <= "10110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111010";
				elsif cntr ="001100111010" THEN
				      t1addb <= "10110011";
				      t2addb <= "10110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111011";
				elsif cntr ="001100111011" THEN
				      t1addb <= "10110100";
				      t2addb <= "10110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111100";
				elsif cntr ="001100111100" THEN
				      t1addb <= "10110101";
				      t2addb <= "10110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111101";
				elsif cntr ="001100111101" THEN
				      t1addb <= "10110110";
				      t2addb <= "10110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111110";
				elsif cntr ="001100111110" THEN
				      t1addb <= "10110111";
				      t2addb <= "10110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001100111111";
				elsif cntr ="001100111111" THEN
				      t1addb <= "10111000";
				      t2addb <= "10111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000000";
				elsif cntr ="001101000000" THEN
				      t1addb <= "10111001";
				      t2addb <= "10111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000001";
				elsif cntr ="001101000001" THEN
				      t1addb <= "10111010";
				      t2addb <= "10111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000010";
				elsif cntr ="001101000010" THEN
				      t1addb <= "10111011";
				      t2addb <= "10111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000011";
				elsif cntr ="001101000011" THEN
				      t1addb <= "10111100";
				      t2addb <= "10111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000100";
				elsif cntr ="001101000100" THEN
				      t1addb <= "10111101";
				      t2addb <= "10111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000101";
				elsif cntr ="001101000101" THEN
				      t1addb <= "10111110";
				      t2addb <= "10111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000110";
				elsif cntr ="001101000110" THEN
				      t1addb <= "10111111";
				      t2addb <= "10111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101000111";
				elsif cntr ="001101000111" THEN
				      t1addb <= "11000000";
				      t2addb <= "11000000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001000";
				elsif cntr ="001101001000" THEN
				      t1addb <= "11000001";
				      t2addb <= "11000001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001001";
				elsif cntr ="001101001001" THEN
				      t1addb <= "11000010";
				      t2addb <= "11000010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001010";
				elsif cntr ="001101001010" THEN
				      t1addb <= "11000011";
				      t2addb <= "11000011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001011";
				elsif cntr ="001101001011" THEN
				      t1addb <= "11000100";
				      t2addb <= "11000100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001100";
				elsif cntr ="001101001100" THEN
				      t1addb <= "11000101";
				      t2addb <= "11000101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001101";
				elsif cntr ="001101001101" THEN
				      t1addb <= "11000110";
				      t2addb <= "11000110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001110";
				elsif cntr ="001101001110" THEN
				      t1addb <= "11000111";
				      t2addb <= "11000111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101001111";
				elsif cntr ="001101001111" THEN
				      t1addb <= "11001000";
				      t2addb <= "11001000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010000";
				elsif cntr ="001101010000" THEN
				      t1addb <= "11001001";
				      t2addb <= "11001001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010001";
				elsif cntr ="001101010001" THEN
				      t1addb <= "11001010";
				      t2addb <= "11001010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010010";
				elsif cntr ="001101010010" THEN
				      t1addb <= "11001011";
				      t2addb <= "11001011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010011";
				elsif cntr ="001101010011" THEN
				      t1addb <= "11001100";
				      t2addb <= "11001100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010100";
				elsif cntr ="001101010100" THEN
				      t1addb <= "11001101";
				      t2addb <= "11001101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010101";
				elsif cntr ="001101010101" THEN
				      t1addb <= "11001110";
				      t2addb <= "11001110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010110";
				elsif cntr ="001101010110" THEN
				      t1addb <= "11001111";
				      t2addb <= "11001111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101010111";
				elsif cntr ="001101010111" THEN
				      t1addb <= "11010000";
				      t2addb <= "11010000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011000";
				elsif cntr ="001101011000" THEN
				      t1addb <= "11010001";
				      t2addb <= "11010001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011001";
				elsif cntr ="001101011001" THEN
				      t1addb <= "11010010";
				      t2addb <= "11010010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011010";
				elsif cntr ="001101011010" THEN
				      t1addb <= "11010011";
				      t2addb <= "11010011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011011";
				elsif cntr ="001101011011" THEN
				      t1addb <= "11010100";
				      t2addb <= "11010100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011100";
				elsif cntr ="001101011100" THEN
				      t1addb <= "11010101";
				      t2addb <= "11010101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011101";
				elsif cntr ="001101011101" THEN
				      t1addb <= "11010110";
				      t2addb <= "11010110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011110";
				elsif cntr ="001101011110" THEN
				      t1addb <= "11010111";
				      t2addb <= "11010111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101011111";
				elsif cntr ="001101011111" THEN
				      t1addb <= "11011000";
				      t2addb <= "11011000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100000";
				elsif cntr ="001101100000" THEN
				      t1addb <= "11011001";
				      t2addb <= "11011001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100001";
				elsif cntr ="001101100001" THEN
				      t1addb <= "11011010";
				      t2addb <= "11011010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100010";
				elsif cntr ="001101100010" THEN
				      t1addb <= "11011011";
				      t2addb <= "11011011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100011";
				elsif cntr ="001101100011" THEN
				      t1addb <= "11011100";
				      t2addb <= "11011100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100100";
				elsif cntr ="001101100100" THEN
				      t1addb <= "11011101";
				      t2addb <= "11011101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100101";
				elsif cntr ="001101100101" THEN
				      t1addb <= "11011110";
				      t2addb <= "11011110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100110";
				elsif cntr ="001101100110" THEN
				      t1addb <= "11011111";
				      t2addb <= "11011111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101100111";
				elsif cntr ="001101100111" THEN
				      t1addb <= "11100000";
				      t2addb <= "11100000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101000";
				elsif cntr ="001101101000" THEN
				      t1addb <= "11100001";
				      t2addb <= "11100001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101001";
				elsif cntr ="001101101001" THEN
				      t1addb <= "11100010";
				      t2addb <= "11100010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101010";
				elsif cntr ="001101101010" THEN
				      t1addb <= "11100011";
				      t2addb <= "11100011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101011";
				elsif cntr ="001101101011" THEN
				      t1addb <= "11100100";
				      t2addb <= "11100100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101100";
				elsif cntr ="001101101100" THEN
				      t1addb <= "11100101";
				      t2addb <= "11100101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101101";
				elsif cntr ="001101101101" THEN
				      t1addb <= "11100110";
				      t2addb <= "11100110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101110";
				elsif cntr ="001101101110" THEN
				      t1addb <= "11100111";
				      t2addb <= "11100111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101101111";
				elsif cntr ="001101101111" THEN
				      t1addb <= "11101000";
				      t2addb <= "11101000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110000";
				elsif cntr ="001101110000" THEN
				      t1addb <= "11101001";
				      t2addb <= "11101001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110001";
				elsif cntr ="001101110001" THEN
				      t1addb <= "11101010";
				      t2addb <= "11101010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110010";
				elsif cntr ="001101110010" THEN
				      t1addb <= "11101011";
				      t2addb <= "11101011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110011";
				elsif cntr ="001101110011" THEN
				      t1addb <= "11101100";
				      t2addb <= "11101100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110100";
				elsif cntr ="001101110100" THEN
				      t1addb <= "11101101";
				      t2addb <= "11101101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110101";
				elsif cntr ="001101110101" THEN
				      t1addb <= "11101110";
				      t2addb <= "11101110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110110";
				elsif cntr ="001101110110" THEN
				      t1addb <= "11101111";
				      t2addb <= "11101111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101110111";
				elsif cntr ="001101110111" THEN
				      t1addb <= "11110000";
				      t2addb <= "11110000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111000";
				elsif cntr ="001101111000" THEN
				      t1addb <= "11110001";
				      t2addb <= "11110001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111001";
				elsif cntr ="001101111001" THEN
				      t1addb <= "11110010";
				      t2addb <= "11110010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111010";
				elsif cntr ="001101111010" THEN
				      t1addb <= "11110011";
				      t2addb <= "11110011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111011";
				elsif cntr ="001101111011" THEN
				      t1addb <= "11110100";
				      t2addb <= "11110100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111100";
				elsif cntr ="001101111100" THEN
				      t1addb <= "11110101";
				      t2addb <= "11110101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111101";
				elsif cntr ="001101111101" THEN
				      t1addb <= "11110110";
				      t2addb <= "11110110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111110";
				elsif cntr ="001101111110" THEN
				      t1addb <= "11110111";
				      t2addb <= "11110111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001101111111";
				elsif cntr ="001101111111" THEN
				      t1addb <= "11111000";
				      t2addb <= "11111000";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000000";
				elsif cntr ="001110000000" THEN
				      t1addb <= "11111001";
				      t2addb <= "11111001";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000001";
				elsif cntr ="001110000001" THEN
				      t1addb <= "11111010";
				      t2addb <= "11111010";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000010";
				elsif cntr ="001110000010" THEN
				      t1addb <= "11111011";
				      t2addb <= "11111011";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000011";
				elsif cntr ="001110000011" THEN
				      t1addb <= "11111100";
				      t2addb <= "11111100";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000100";
				elsif cntr ="001110000100" THEN
				      t1addb <= "11111101";
				      t2addb <= "11111101";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000101";
				elsif cntr ="001110000101" THEN
				      t1addb <= "11111110";
				      t2addb <= "11111110";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000110";
				elsif cntr ="001110000110" THEN
				      t1addb <= "11111111";
				      t2addb <= "11111111";
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110000111";
				elsif cntr ="001110000111" THEN
				      
				      
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001000";
				elsif cntr ="001110001000" THEN
				      
				      
				      bfrjin   <= t1doutb;
				      bfrjplin <= t2doutb;
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001001";
				elsif cntr ="001110001001" THEN
				      
				      
				      
				      
				      
				      
				      
				      
				      
				      
				      cntr <= "001110001010";
				elsif cntr ="001110001010" THEN
				      
				      
				   
				   
				   
				   
				   
				   
				   
				   
				   
				      
				      
				      
				      cntr <= "001110001011";
				elsif cntr ="001110001011" THEN
				
					
					
					
				     pdone <= '1';
				   
				   
				   
					
					 cntr <= "001110001100";
				elsif cntr ="001110001100" THEN
				
				
					cntr <= "000000000000";
				
				






				END IF;
				
				
				
								
				if cntr1 ="000000000000" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000001" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000010" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000011" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000100" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000101" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000110" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000000111" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="000000001000" THEN
				
				
				
					  t1wea <= '1';
				      
				      t1adda <= "00000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000000111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001000111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000001111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010000010" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111010";
				      
				      
				      t1dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="000010000011" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111011";
				      
				      
				      t1dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="000010000100" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111100";
				      
				      
				      t1dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="000010000101" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111101";
				      
				      
				      t1dina <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="000010000110" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111110";
				      
				      
				      t1dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000010000111" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111111";
				      
				      
				      t1dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000010001000" THEN
				
				
				
					  t2wea <= '1';
				      
				      t2adda <= "00000000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010001111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00000111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010010111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00001111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010011111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00010111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010100111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00011111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010101111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00100111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010110111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00101111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000010111111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00110111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011000111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "00111111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011001111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01000111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011010111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01001111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011011111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01010111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011100111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01011111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011101111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01100111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011110111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01101111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000011111111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01110111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100000000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100000001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100000010" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111010";
				      
				      
				      t2dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="000100000011" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111011";
				      
				      
				      t2dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="000100000100" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111100";
				      
				      
				      t2dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="000100000101" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111101";
				      
				      
				      t2dina <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="000100000110" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111110";
				      
				      
				      t2dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000100000111" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "01111111";
				      
				      
				      t2dina <= bfrjplout;
				                                   
				                                   
				                                   
				elsif cntr1 ="000100001000" THEN
				
				
				
					  t1wea <= '1';
				      
				      t1adda <= "10000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000100111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101000111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "10111111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000101111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110000010" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111010";
				      
				      
				      t1dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="000110000011" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111011";
				      
				      
				      t1dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="000110000100" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111100";
				      
				      
				      t1dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="000110000101" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111101";
				      
				      
				      t1dina <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="000110000110" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111110";
				      
				      
				      t1dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="000110000111" THEN 
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "11111111";
				      
				      
				      t1dina <= bfrjplout;
				                                   
				                                   
				                                   
				elsif cntr1 ="000110001000" THEN
				
				
				
					  t2wea <= '1';
				      
				      t2adda <= "10000000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110001111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10000111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110010111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10001111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110011111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10010111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110100111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10011111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110101111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10100111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110110111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10101111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000110111111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10110111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111000111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "10111111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111001111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11000111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111010111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11001111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111011111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11010111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111100111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11011111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111101111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11100111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111110111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11101111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111010" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110010";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111011" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110011";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111100" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110100";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111101" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110101";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111110" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110110";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="000111111111" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11110111";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000000000" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111000";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000000001" THEN
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111001";
				      
				      
				      t2dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000000010" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111010";
				      
				      
				      t2dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="001000000011" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111011";
				      
				      
				      t2dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="001000000100" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111100";
				      
				      
				      t2dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="001000000101" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111101";
				      
				      
				      t2dina <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="001000000110" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111110";
				      
				      
				      t2dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001000000111" THEN 
				      
				      
				      
				      t2wea <= '1';
				      
				      t2adda <= "11111111";
				      
				      
				      t2dina <= bfrjplout;
				                                  
				                                  
				                                  
				elsif cntr1 ="001000001000" THEN
				
				
				
					  t1wea <= '1';
				      
				      t1adda <= "00000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001000111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001000111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "00111111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001001111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01000111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001010111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01001111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001011111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01010111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001100111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01011111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001101111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01100111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001110111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01101111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110010";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110011";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110100";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110101";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110110";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001001111111" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01110111";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010000000" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111000";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010000001" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111001";
				      
				      
				      t1dina <= bfrjplout;
				      
				      
				      
				elsif cntr1 ="001010000010" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111010";
				      
				      
				      t1dina <= bfrjplout;
				            
				            
				            
				elsif cntr1 ="001010000011" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111011";
				      
				      
				      t1dina <= bfrjplout;
				                  
				                  
				                  
				elsif cntr1 ="001010000100" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111100";
				      
				      
				      t1dina <= bfrjplout;
				                        
				                        
				                        
				elsif cntr1 ="001010000101" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111101";
				      
				      
				      t1dina <= bfrjplout;
				                              
				                              
				                              
				elsif cntr1 ="001010000110" THEN
				      
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111110";
				      
				      
				      t1dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001010000111" THEN
				      
				      
				      t1wea <= '1';
				      
				      t1adda <= "01111111";
				      
				      
				      t1dina <= bfrjplout;
				                                    
				                                    
				                                    
				elsif cntr1 ="001010001000" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="001010001001" THEN
				
				
				
				
				
				
				
				
				
				
				
				
				elsif cntr1 ="001010001010" THEN
				
				
				
					  ioweb <= '1';
				      
				      ioaddb <= "000000000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001010111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011000111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001011111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111000";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100000111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111010";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111100";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001001" THEN 
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111110";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001010" THEN
				
				
				
					  ioweb <= '1';
				      
				      ioaddb <= "000000001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000000111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000001111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000010111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000011111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000100111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000101111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000110111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "000111111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001000111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001001111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001010111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001011111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001100111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001100111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001101111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001110111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101000111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "001111111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010000111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101001111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010001111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010010111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101010111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010011111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010100111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101011111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010101111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010110111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101100111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "010111111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011000111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101101111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011001111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011010111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101110111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011011111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011100111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001101111111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011101111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000010" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000011" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000100" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000101" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011110111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000110" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111001";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110000111" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111011";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110001000" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111101";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110001001" THEN
				      
				      
				      
				      ioweb <= '1';
				      
				      ioaddb <= "011111111";
				      
				      
				      iodinb <= bfrjout;
				      
				      
				      
				elsif cntr1 ="001110001010" THEN
				   
				   
				   
		
		



				   
				      
				      
				      
				elsif cntr1 ="001110001011" THEN
				
				









				
				END IF;
				











			
				
				
				
				
				
				
				
			
			END IF;
			
		
		
		END IF;
	
	
  END IF;	
 
 
END PROCESS;







 PROCESS (cur_st, en, pdone , mode )
  BEGIN
   
   nxt_st <= cur_st;
   
   done<='0';
   
   busy<='1';

   
    CASE cur_st  IS
      WHEN idle =>
		
		busy<='0';
		

		
		IF en = '1'   THEN
		
			IF mode	="00" THEN
		
				nxt_st <= tontt;
		
			END IF;
			
			IF mode	="10" THEN
			
				nxt_st <= toinvntt;
			
			END IF;
			
			IF mode	="01" THEN
			
				nxt_st <= topwm;
			
			END IF;
		
		END IF;
		
		

	  
	  
      WHEN tontt =>
			
			
			IF pdone = '1'   THEN
		
			nxt_st <= idle;
			
			done <='1';
		
			END IF;

			
      WHEN toinvntt =>
		

		
			IF pdone = '1'   THEN
		
			nxt_st <= idle;
			
			done <='1';
		
			END IF;
			
			
			
			
	  WHEN topwm =>

		
			IF pdone = '1'   THEN
		
			nxt_st <= idle;
			
			done <='1';
		
			END IF;
			
	  
	
		
    END CASE;  
	
END PROCESS;
	












 
 END behaviour;